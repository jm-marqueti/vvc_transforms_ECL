module dst7_8(
input signed [8:0]X[7:0],
output signed [15:0]Y[7:0]);

// SAU
/*

// Adder Trees
assign Y[0] = x11[0] + x22[1] + x33[2] + x42[3] + x50[4] + x56[5] + x60[6] + x62[7];
assign Y[1] = x33[0] + x56[1] + x62[2] + x50[3] + x22[4] - x11[5] - x42[6] - x60[7];
assign Y[2] = x50[0] + x60[1] + x22[2] - x33[3] - x62[4] - x42[5] + x11[6] + x56[7];
assign Y[3] = x60[0] + x33[1] - x42[2] - x56[3] + x11[4] + x62[5] + x22[6] - x50[7];
assign Y[4] = x62[0] - x11[1] - x60[2] + x22[3] + x56[4] - x33[5] - x50[6] + x42[7];
assign Y[5] = x56[0] - x50[1] - x11[2] + x60[3] - x42[4] - x22[5] + x62[6] - x33[7];
assign Y[6] = x42[0] - x62[1] + x50[2] - x11[3] - x33[4] + x60[5] - x56[6] + x22[7];
assign Y[7] = x22[0] - x42[1] + x56[2] - x62[3] + x60[4] - x50[5] + x33[6] - x11[7];

*/

endmodule