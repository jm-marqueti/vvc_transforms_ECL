module decomp_1 (input signed [16:0]a,b,
output signed [17:0] even, odd);

assign even = a + b;

assign odd = a - b;

endmodule