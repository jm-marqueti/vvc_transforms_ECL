module dst7_1d(
input [8:0]X[31:0],
input [1:0]N,
output [15:0]Y[31:0]);




endmodule