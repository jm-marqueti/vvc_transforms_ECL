module dst7_32(
input signed [8:0]X[31:0],
output signed [15:0]Y[31:0]);

// SAU
/*
// Adder Trees
assign Y[0] = x2[0] + x3[1] + x5[2] + x6[3] + x8[4] + x9[5] + x11[6] + x12[7] + x13[8] + x15[9] + x16[10] + x17[11] + x19[12] + x20[13] + x21[14] + x22[15] + x23[16] + x24[17] + x25[18] + x26[19] + x27[20] + x28[21] + x28[22] + x29[23] + x30[24] + x30[25] + x31[26] + x31[27] + x31[28] + x32[29] + x32[30] + x32[31];
assign Y[1] = x5[0] + x9[1] + x13[2] + x17[3] + x21[4] + x24[5] + x27[6] + x29[7] + x31[8] + x32[9] + x32[10] + x31[11] + x30[12] + x28[13] + x26[14] + x23[15] + x20[16] + x16[17] + x12[18] + x8[19] + x3[20] - x2[21] - x6[22] - x11[23] - x15[24] - x19[25] - x22[26] - x25[27] - x28[28] - x30[29] - x31[30] - x32[31];
assign Y[2] = x8[0] + x15[1] + x21[2] + x26[3] + x30[4] + x32[5] + x32[6] + x30[7] + x26[8] + x21[9] + x15[10] + x8[11] - x8[13] - x15[14] - x21[15] - x26[16] - x30[17] - x32[18] - x32[19] - x30[20] - x26[21] - x21[22] - x15[23] - x8[24] + x8[26] + x15[27] + x21[28] + x26[29] + x30[30] + x32[31];
assign Y[3] = x11[0] + x20[1] + x27[2] + x31[3] + x32[4] + x28[5] + x22[6] + x13[7] + x3[8] - x8[9] - x17[10] - x25[11] - x30[12] - x32[13] - x30[14] - x24[15] - x16[16] - x6[17] + x5[18] + x15[19] + x23[20] + x29[21] + x32[22] + x31[23] + x26[24] + x19[25] + x9[26] - x2[27] - x12[28] - x21[29] - x28[30] - x31[31];
assign Y[4] = x13[0] + x24[1] + x31[2] + x31[3] + x26[4] + x16[5] + x3[6] - x11[7] - x22[8] - x30[9] - x32[10] - x28[11] - x19[12] - x6[13] + x8[14] + x20[15] + x28[16] + x32[17] + x29[18] + x21[19] + x9[20] - x5[21] - x17[22] - x27[23] - x32[24] - x30[25] - x23[26] - x12[27] + x2[28] + x15[29] + x25[30] + x31[31];
assign Y[5] = x16[0] + x28[1] + x32[2] + x27[3] + x15[4] - x2[5] - x17[6] - x28[7] - x32[8] - x26[9] - x13[10] + x3[11] + x19[12] + x29[13] + x32[14] + x25[15] + x12[16] - x5[17] - x20[18] - x30[19] - x31[20] - x24[21] - x11[22] + x6[23] + x21[24] + x30[25] + x31[26] + x23[27] + x9[28] - x8[29] - x22[30] - x31[31];
assign Y[6] = x19[0] + x30[1] + x30[2] + x19[3] - x19[5] - x30[6] - x30[7] - x19[8] + x19[10] + x30[11] + x30[12] + x19[13] - x19[15] - x30[16] - x30[17] - x19[18] + x19[20] + x30[21] + x30[22] + x19[23] - x19[25] - x30[26] - x30[27] - x19[28] + x19[30] + x30[31];
assign Y[7] = x21[0] + x32[1] + x26[2] + x8[3] - x15[4] - x30[5] - x30[6] - x15[7] + x8[8] + x26[9] + x32[10] + x21[11] - x21[13] - x32[14] - x26[15] - x8[16] + x15[17] + x30[18] + x30[19] + x15[20] - x8[21] - x26[22] - x32[23] - x21[24] + x21[26] + x32[27] + x26[28] + x8[29] - x15[30] - x30[31];
assign Y[8] = x23[0] + x32[1] + x20[2] - x5[3] - x26[4] - x31[5] - x16[6] + x9[7] + x28[8] + x30[9] + x12[10] - x13[11] - x30[12] - x28[13] - x8[14] + x17[15] + x31[16] + x25[17] + x3[18] - x21[19] - x32[20] - x22[21] + x2[22] + x24[23] + x32[24] + x19[25] - x6[26] - x27[27] - x31[28] - x15[29] + x11[30] + x29[31];
assign Y[9] = x25[0] + x31[1] + x12[2] - x16[3] - x32[4] - x22[5] + x5[6] + x28[7] + x29[8] + x8[9] - x20[10] - x32[11] - x19[12] + x9[13] + x30[14] + x27[15] + x3[16] - x23[17] - x31[18] - x15[19] + x13[20] + x31[21] + x24[22] - x2[23] - x26[24] - x30[25] - x11[26] + x17[27] + x32[28] + x21[29] - x6[30] - x28[31];
assign Y[10] = x27[0] + x28[1] + x3[2] - x25[3] - x30[4] - x6[5] + x23[6] + x31[7] + x9[8] - x21[9] - x31[10] - x12[11] + x19[12] + x32[13] + x15[14] - x16[15] - x32[16] - x17[17] + x13[18] + x32[19] + x20[20] - x11[21] - x31[22] - x22[23] + x8[24] + x30[25] + x24[26] - x5[27] - x29[28] - x26[29] + x2[30] + x28[31];
assign Y[11] = x28[0] + x25[1] - x6[2] - x31[3] - x21[4] + x12[5] + x32[6] + x16[7] - x17[8] - x32[9] - x11[10] + x22[11] + x30[12] + x5[13] - x26[14] - x28[15] + x2[16] + x29[17] + x24[18] - x8[19] - x31[20] - x20[21] + x13[22] + x32[23] + x15[24] - x19[25] - x31[26] - x9[27] + x23[28] + x30[29] + x3[30] - x27[31];
assign Y[12] = x30[0] + x21[1] - x15[2] - x32[3] - x8[4] + x26[5] + x26[6] - x8[7] - x32[8] - x15[9] + x21[10] + x30[11] - x30[13] - x21[14] + x15[15] + x32[16] + x8[17] - x26[18] - x26[19] + x8[20] + x32[21] + x15[22] - x21[23] - x30[24] + x30[26] + x21[27] - x15[28] - x32[29] - x8[30] + x26[31];
assign Y[13] = x31[0] + x16[1] - x22[2] - x28[3] + x8[4] + x32[5] + x9[6] - x27[7] - x23[8] + x15[9] + x31[10] + x2[11] - x30[12] - x17[13] + x21[14] + x28[15] - x6[16] - x32[17] - x11[18] + x26[19] + x24[20] - x13[21] - x31[22] - x3[23] + x30[24] + x19[25] - x20[26] - x29[27] + x5[28] + x32[29] + x12[30] - x25[31];
assign Y[14] = x31[0] + x11[1] - x28[2] - x20[3] + x21[4] + x27[5] - x12[6] - x31[7] + x2[8] + x32[9] + x9[10] - x28[11] - x19[12] + x22[13] + x26[14] - x13[15] - x31[16] + x3[17] + x32[18] + x8[19] - x29[20] - x17[21] + x23[22] + x25[23] - x15[24] - x30[25] + x5[26] + x32[27] + x6[28] - x30[29] - x16[30] + x24[31];
assign Y[15] = x32[0] + x5[1] - x31[2] - x9[3] + x30[4] + x13[5] - x28[6] - x17[7] + x25[8] + x21[9] - x22[10] - x24[11] + x19[12] + x27[13] - x15[14] - x29[15] + x11[16] + x31[17] - x6[18] - x32[19] + x2[20] + x32[21] + x3[22] - x31[23] - x8[24] + x30[25] + x12[26] - x28[27] - x16[28] + x26[29] + x20[30] - x23[31];
assign Y[16] = x32[0] - x2[1] - x32[2] + x3[3] + x32[4] - x5[5] - x31[6] + x6[7] + x31[8] - x8[9] - x31[10] + x9[11] + x30[12] - x11[13] - x30[14] + x12[15] + x29[16] - x13[17] - x28[18] + x15[19] + x28[20] - x16[21] - x27[22] + x17[23] + x26[24] - x19[25] - x25[26] + x20[27] + x24[28] - x21[29] - x23[30] + x22[31];
assign Y[17] = x32[0] - x8[1] - x30[2] + x15[3] + x26[4] - x21[5] - x21[6] + x26[7] + x15[8] - x30[9] - x8[10] + x32[11] - x32[13] + x8[14] + x30[15] - x15[16] - x26[17] + x21[18] + x21[19] - x26[20] - x15[21] + x30[22] + x8[23] - x32[24] + x32[26] - x8[27] - x30[28] + x15[29] + x26[30] - x21[31];
assign Y[18] = x31[0] - x13[1] - x25[2] + x24[3] + x15[4] - x31[5] - x2[6] + x31[7] - x12[8] - x26[9] + x23[10] + x16[11] - x30[12] - x3[13] + x32[14] - x11[15] - x27[16] + x22[17] + x17[18] - x30[19] - x5[20] + x32[21] - x9[22] - x28[23] + x21[24] + x19[25] - x29[26] - x6[27] + x32[28] - x8[29] - x28[30] + x20[31];
assign Y[19] = x30[0] - x19[1] - x19[2] + x30[3] - x30[5] + x19[6] + x19[7] - x30[8] + x30[10] - x19[11] - x19[12] + x30[13] - x30[15] + x19[16] + x19[17] - x30[18] + x30[20] - x19[21] - x19[22] + x30[23] - x30[25] + x19[26] + x19[27] - x30[28] + x30[30] - x19[31];
assign Y[20] = x29[0] - x23[1] - x11[2] + x32[3] - x15[4] - x20[5] + x31[6] - x5[7] - x27[8] + x26[9] + x6[10] - x31[11] + x19[12] + x16[13] - x32[14] + x9[15] + x24[16] - x28[17] - x2[18] + x30[19] - x22[20] - x12[21] + x32[22] - x13[23] - x21[24] + x30[25] - x3[26] - x28[27] + x25[28] + x8[29] - x31[30] + x17[31];
assign Y[21] = x28[0] - x27[1] - x2[2] + x28[3] - x26[4] - x3[5] + x29[6] - x25[7] - x5[8] + x30[9] - x24[10] - x6[11] + x30[12] - x23[13] - x8[14] + x31[15] - x22[16] - x9[17] + x31[18] - x21[19] - x11[20] + x31[21] - x20[22] - x12[23] + x32[24] - x19[25] - x13[26] + x32[27] - x17[28] - x15[29] + x32[30] - x16[31];
assign Y[22] = x26[0] - x30[1] + x8[2] + x21[3] - x32[4] + x15[5] + x15[6] - x32[7] + x21[8] + x8[9] - x30[10] + x26[11] - x26[13] + x30[14] - x8[15] - x21[16] + x32[17] - x15[18] - x15[19] + x32[20] - x21[21] - x8[22] + x30[23] - x26[24] + x26[26] - x30[27] + x8[28] + x21[29] - x32[30] + x15[31];
assign Y[23] = x24[0] - x31[1] + x16[2] + x11[3] - x30[4] + x28[5] - x6[6] - x20[7] + x32[8] - x21[9] - x5[10] + x27[11] - x30[12] + x12[13] + x15[14] - x31[15] + x25[16] - x2[17] - x23[18] + x32[19] - x17[20] - x9[21] + x29[22] - x28[23] + x8[24] + x19[25] - x32[26] + x22[27] + x3[28] - x26[29] + x31[30] - x13[31];
assign Y[24] = x22[0] - x32[1] + x23[2] - x2[3] - x21[4] + x32[5] - x24[6] + x3[7] + x20[8] - x32[9] + x25[10] - x5[11] - x19[12] + x31[13] - x26[14] + x6[15] + x17[16] - x31[17] + x27[18] - x8[19] - x16[20] + x31[21] - x28[22] + x9[23] + x15[24] - x30[25] + x28[26] - x11[27] - x13[28] + x30[29] - x29[30] + x12[31];
assign Y[25] = x20[0] - x31[1] + x28[2] - x13[3] - x8[4] + x25[5] - x32[6] + x24[7] - x6[8] - x15[9] + x29[10] - x31[11] + x19[12] + x2[13] - x21[14] + x31[15] - x28[16] + x12[17] + x9[18] - x26[19] + x32[20] - x23[21] + x5[22] + x16[23] - x30[24] + x30[25] - x17[26] - x3[27] + x22[28] - x32[29] + x27[30] - x11[31];
assign Y[26] = x17[0] - x29[1] + x31[2] - x23[3] + x8[4] + x11[5] - x25[6] + x32[7] - x28[8] + x15[9] + x3[10] - x20[11] + x30[12] - x31[13] + x21[14] - x5[15] - x13[16] + x27[17] - x32[18] + x26[19] - x12[20] - x6[21] + x22[22] - x31[23] + x30[24] - x19[25] + x2[26] + x16[27] - x28[28] + x32[29] - x24[30] + x9[31];
assign Y[27] = x15[0] - x26[1] + x32[2] - x30[3] + x21[4] - x8[5] - x8[6] + x21[7] - x30[8] + x32[9] - x26[10] + x15[11] - x15[13] + x26[14] - x32[15] + x30[16] - x21[17] + x8[18] + x8[19] - x21[20] + x30[21] - x32[22] + x26[23] - x15[24] + x15[26] - x26[27] + x32[28] - x30[29] + x21[30] - x8[31];
assign Y[28] = x12[0] - x22[1] + x29[2] - x32[3] + x30[4] - x23[5] + x13[6] - x2[7] - x11[8] + x21[9] - x28[10] + x32[11] - x30[12] + x24[13] - x15[14] + x3[15] + x9[16] - x20[17] + x28[18] - x32[19] + x31[20] - x25[21] + x16[22] - x5[23] - x8[24] + x19[25] - x27[26] + x31[27] - x31[28] + x26[29] - x17[30] + x6[31];
assign Y[29] = x9[0] - x17[1] + x24[2] - x29[3] + x32[4] - x31[5] + x28[6] - x23[7] + x16[8] - x8[9] - x2[10] + x11[11] - x19[12] + x25[13] - x30[14] + x32[15] - x31[16] + x28[17] - x22[18] + x15[19] - x6[20] - x3[21] + x12[22] - x20[23] + x26[24] - x30[25] + x32[26] - x31[27] + x27[28] - x21[29] + x13[30] - x5[31];
assign Y[30] = x6[0] - x12[1] + x17[2] - x22[3] + x26[4] - x29[5] + x31[6] - x32[7] + x31[8] - x30[9] + x27[10] - x23[11] + x19[12] - x13[13] + x8[14] - x2[15] - x5[16] + x11[17] - x16[18] + x21[19] - x25[20] + x28[21] - x31[22] + x32[23] - x32[24] + x30[25] - x28[26] + x24[27] - x20[28] + x15[29] - x9[30] + x3[31];
assign Y[31] = x3[0] - x6[1] + x9[2] - x12[3] + x15[4] - x17[5] + x20[6] - x22[7] + x24[8] - x26[9] + x28[10] - x29[11] + x30[12] - x31[13] + x32[14] - x32[15] + x32[16] - x31[17] + x31[18] - x30[19] + x28[20] - x27[21] + x25[22] - x23[23] + x21[24] - x19[25] + x16[26] - x13[27] + x11[28] - x8[29] + x5[30] - x2[31];

*/
endmodule