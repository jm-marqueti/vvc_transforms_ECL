module transpose_buffer_32x32 (
	clock, 
	reset,
	enable,
	direction,
	in_buffer,
	out_0,
	out_1,
	out_2,
	out_3,
	out_4,
	out_5,
	out_6,
	out_7,
	out_8,
	out_9,
	out_10,
	out_11,
	out_12,
	out_13,
	out_14,
	out_15,
	out_16,
	out_17,
	out_18,
	out_19,
	out_20,
	out_21,
	out_22,
	out_23,
	out_24,
	out_25,
	out_26,
	out_27,
	out_28,
	out_29,
	out_30,
	out_31
);

parameter DATA_WIDTH = 16;
input  clock, reset, enable, direction;
input  [(32*DATA_WIDTH)-1:0] in_buffer;
wire  [DATA_WIDTH-1:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27, in_28, in_29, in_30, in_31;
output [DATA_WIDTH-1:0] out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, out_11, out_12, out_13, out_14, out_15, out_16, out_17, out_18, out_19, out_20, out_21, out_22, out_23, out_24, out_25, out_26, out_27, out_28, out_29, out_30, out_31;
wire   [DATA_WIDTH-1:0] out_of_0_0, out_of_0_1, out_of_0_2, out_of_0_3, out_of_0_4, out_of_0_5, out_of_0_6, out_of_0_7, out_of_0_8, out_of_0_9, out_of_0_10, out_of_0_11, out_of_0_12, out_of_0_13, out_of_0_14, out_of_0_15, out_of_0_16, out_of_0_17, out_of_0_18, out_of_0_19, out_of_0_20, out_of_0_21, out_of_0_22, out_of_0_23, out_of_0_24, out_of_0_25, out_of_0_26, out_of_0_27, out_of_0_28, out_of_0_29, out_of_0_30, out_of_0_31, out_of_1_0, out_of_1_1, out_of_1_2, out_of_1_3, out_of_1_4, out_of_1_5, out_of_1_6, out_of_1_7, out_of_1_8, out_of_1_9, out_of_1_10, out_of_1_11, out_of_1_12, out_of_1_13, out_of_1_14, out_of_1_15, out_of_1_16, out_of_1_17, out_of_1_18, out_of_1_19, out_of_1_20, out_of_1_21, out_of_1_22, out_of_1_23, out_of_1_24, out_of_1_25, out_of_1_26, out_of_1_27, out_of_1_28, out_of_1_29, out_of_1_30, out_of_1_31, out_of_2_0, out_of_2_1, out_of_2_2, out_of_2_3, out_of_2_4, out_of_2_5, out_of_2_6, out_of_2_7, out_of_2_8, out_of_2_9, out_of_2_10, out_of_2_11, out_of_2_12, out_of_2_13, out_of_2_14, out_of_2_15, out_of_2_16, out_of_2_17, out_of_2_18, out_of_2_19, out_of_2_20, out_of_2_21, out_of_2_22, out_of_2_23, out_of_2_24, out_of_2_25, out_of_2_26, out_of_2_27, out_of_2_28, out_of_2_29, out_of_2_30, out_of_2_31, out_of_3_0, out_of_3_1, out_of_3_2, out_of_3_3, out_of_3_4, out_of_3_5, out_of_3_6, out_of_3_7, out_of_3_8, out_of_3_9, out_of_3_10, out_of_3_11, out_of_3_12, out_of_3_13, out_of_3_14, out_of_3_15, out_of_3_16, out_of_3_17, out_of_3_18, out_of_3_19, out_of_3_20, out_of_3_21, out_of_3_22, out_of_3_23, out_of_3_24, out_of_3_25, out_of_3_26, out_of_3_27, out_of_3_28, out_of_3_29, out_of_3_30, out_of_3_31, out_of_4_0, out_of_4_1, out_of_4_2, out_of_4_3, out_of_4_4, out_of_4_5, out_of_4_6, out_of_4_7, out_of_4_8, out_of_4_9, out_of_4_10, out_of_4_11, out_of_4_12, out_of_4_13, out_of_4_14, out_of_4_15, out_of_4_16, out_of_4_17, out_of_4_18, out_of_4_19, out_of_4_20, out_of_4_21, out_of_4_22, out_of_4_23, out_of_4_24, out_of_4_25, out_of_4_26, out_of_4_27, out_of_4_28, out_of_4_29, out_of_4_30, out_of_4_31, out_of_5_0, out_of_5_1, out_of_5_2, out_of_5_3, out_of_5_4, out_of_5_5, out_of_5_6, out_of_5_7, out_of_5_8, out_of_5_9, out_of_5_10, out_of_5_11, out_of_5_12, out_of_5_13, out_of_5_14, out_of_5_15, out_of_5_16, out_of_5_17, out_of_5_18, out_of_5_19, out_of_5_20, out_of_5_21, out_of_5_22, out_of_5_23, out_of_5_24, out_of_5_25, out_of_5_26, out_of_5_27, out_of_5_28, out_of_5_29, out_of_5_30, out_of_5_31, out_of_6_0, out_of_6_1, out_of_6_2, out_of_6_3, out_of_6_4, out_of_6_5, out_of_6_6, out_of_6_7, out_of_6_8, out_of_6_9, out_of_6_10, out_of_6_11, out_of_6_12, out_of_6_13, out_of_6_14, out_of_6_15, out_of_6_16, out_of_6_17, out_of_6_18, out_of_6_19, out_of_6_20, out_of_6_21, out_of_6_22, out_of_6_23, out_of_6_24, out_of_6_25, out_of_6_26, out_of_6_27, out_of_6_28, out_of_6_29, out_of_6_30, out_of_6_31, out_of_7_0, out_of_7_1, out_of_7_2, out_of_7_3, out_of_7_4, out_of_7_5, out_of_7_6, out_of_7_7, out_of_7_8, out_of_7_9, out_of_7_10, out_of_7_11, out_of_7_12, out_of_7_13, out_of_7_14, out_of_7_15, out_of_7_16, out_of_7_17, out_of_7_18, out_of_7_19, out_of_7_20, out_of_7_21, out_of_7_22, out_of_7_23, out_of_7_24, out_of_7_25, out_of_7_26, out_of_7_27, out_of_7_28, out_of_7_29, out_of_7_30, out_of_7_31, out_of_8_0, out_of_8_1, out_of_8_2, out_of_8_3, out_of_8_4, out_of_8_5, out_of_8_6, out_of_8_7, out_of_8_8, out_of_8_9, out_of_8_10, out_of_8_11, out_of_8_12, out_of_8_13, out_of_8_14, out_of_8_15, out_of_8_16, out_of_8_17, out_of_8_18, out_of_8_19, out_of_8_20, out_of_8_21, out_of_8_22, out_of_8_23, out_of_8_24, out_of_8_25, out_of_8_26, out_of_8_27, out_of_8_28, out_of_8_29, out_of_8_30, out_of_8_31, out_of_9_0, out_of_9_1, out_of_9_2, out_of_9_3, out_of_9_4, out_of_9_5, out_of_9_6, out_of_9_7, out_of_9_8, out_of_9_9, out_of_9_10, out_of_9_11, out_of_9_12, out_of_9_13, out_of_9_14, out_of_9_15, out_of_9_16, out_of_9_17, out_of_9_18, out_of_9_19, out_of_9_20, out_of_9_21, out_of_9_22, out_of_9_23, out_of_9_24, out_of_9_25, out_of_9_26, out_of_9_27, out_of_9_28, out_of_9_29, out_of_9_30, out_of_9_31, out_of_10_0, out_of_10_1, out_of_10_2, out_of_10_3, out_of_10_4, out_of_10_5, out_of_10_6, out_of_10_7, out_of_10_8, out_of_10_9, out_of_10_10, out_of_10_11, out_of_10_12, out_of_10_13, out_of_10_14, out_of_10_15, out_of_10_16, out_of_10_17, out_of_10_18, out_of_10_19, out_of_10_20, out_of_10_21, out_of_10_22, out_of_10_23, out_of_10_24, out_of_10_25, out_of_10_26, out_of_10_27, out_of_10_28, out_of_10_29, out_of_10_30, out_of_10_31, out_of_11_0, out_of_11_1, out_of_11_2, out_of_11_3, out_of_11_4, out_of_11_5, out_of_11_6, out_of_11_7, out_of_11_8, out_of_11_9, out_of_11_10, out_of_11_11, out_of_11_12, out_of_11_13, out_of_11_14, out_of_11_15, out_of_11_16, out_of_11_17, out_of_11_18, out_of_11_19, out_of_11_20, out_of_11_21, out_of_11_22, out_of_11_23, out_of_11_24, out_of_11_25, out_of_11_26, out_of_11_27, out_of_11_28, out_of_11_29, out_of_11_30, out_of_11_31, out_of_12_0, out_of_12_1, out_of_12_2, out_of_12_3, out_of_12_4, out_of_12_5, out_of_12_6, out_of_12_7, out_of_12_8, out_of_12_9, out_of_12_10, out_of_12_11, out_of_12_12, out_of_12_13, out_of_12_14, out_of_12_15, out_of_12_16, out_of_12_17, out_of_12_18, out_of_12_19, out_of_12_20, out_of_12_21, out_of_12_22, out_of_12_23, out_of_12_24, out_of_12_25, out_of_12_26, out_of_12_27, out_of_12_28, out_of_12_29, out_of_12_30, out_of_12_31, out_of_13_0, out_of_13_1, out_of_13_2, out_of_13_3, out_of_13_4, out_of_13_5, out_of_13_6, out_of_13_7, out_of_13_8, out_of_13_9, out_of_13_10, out_of_13_11, out_of_13_12, out_of_13_13, out_of_13_14, out_of_13_15, out_of_13_16, out_of_13_17, out_of_13_18, out_of_13_19, out_of_13_20, out_of_13_21, out_of_13_22, out_of_13_23, out_of_13_24, out_of_13_25, out_of_13_26, out_of_13_27, out_of_13_28, out_of_13_29, out_of_13_30, out_of_13_31, out_of_14_0, out_of_14_1, out_of_14_2, out_of_14_3, out_of_14_4, out_of_14_5, out_of_14_6, out_of_14_7, out_of_14_8, out_of_14_9, out_of_14_10, out_of_14_11, out_of_14_12, out_of_14_13, out_of_14_14, out_of_14_15, out_of_14_16, out_of_14_17, out_of_14_18, out_of_14_19, out_of_14_20, out_of_14_21, out_of_14_22, out_of_14_23, out_of_14_24, out_of_14_25, out_of_14_26, out_of_14_27, out_of_14_28, out_of_14_29, out_of_14_30, out_of_14_31, out_of_15_0, out_of_15_1, out_of_15_2, out_of_15_3, out_of_15_4, out_of_15_5, out_of_15_6, out_of_15_7, out_of_15_8, out_of_15_9, out_of_15_10, out_of_15_11, out_of_15_12, out_of_15_13, out_of_15_14, out_of_15_15, out_of_15_16, out_of_15_17, out_of_15_18, out_of_15_19, out_of_15_20, out_of_15_21, out_of_15_22, out_of_15_23, out_of_15_24, out_of_15_25, out_of_15_26, out_of_15_27, out_of_15_28, out_of_15_29, out_of_15_30, out_of_15_31, out_of_16_0, out_of_16_1, out_of_16_2, out_of_16_3, out_of_16_4, out_of_16_5, out_of_16_6, out_of_16_7, out_of_16_8, out_of_16_9, out_of_16_10, out_of_16_11, out_of_16_12, out_of_16_13, out_of_16_14, out_of_16_15, out_of_16_16, out_of_16_17, out_of_16_18, out_of_16_19, out_of_16_20, out_of_16_21, out_of_16_22, out_of_16_23, out_of_16_24, out_of_16_25, out_of_16_26, out_of_16_27, out_of_16_28, out_of_16_29, out_of_16_30, out_of_16_31, out_of_17_0, out_of_17_1, out_of_17_2, out_of_17_3, out_of_17_4, out_of_17_5, out_of_17_6, out_of_17_7, out_of_17_8, out_of_17_9, out_of_17_10, out_of_17_11, out_of_17_12, out_of_17_13, out_of_17_14, out_of_17_15, out_of_17_16, out_of_17_17, out_of_17_18, out_of_17_19, out_of_17_20, out_of_17_21, out_of_17_22, out_of_17_23, out_of_17_24, out_of_17_25, out_of_17_26, out_of_17_27, out_of_17_28, out_of_17_29, out_of_17_30, out_of_17_31, out_of_18_0, out_of_18_1, out_of_18_2, out_of_18_3, out_of_18_4, out_of_18_5, out_of_18_6, out_of_18_7, out_of_18_8, out_of_18_9, out_of_18_10, out_of_18_11, out_of_18_12, out_of_18_13, out_of_18_14, out_of_18_15, out_of_18_16, out_of_18_17, out_of_18_18, out_of_18_19, out_of_18_20, out_of_18_21, out_of_18_22, out_of_18_23, out_of_18_24, out_of_18_25, out_of_18_26, out_of_18_27, out_of_18_28, out_of_18_29, out_of_18_30, out_of_18_31, out_of_19_0, out_of_19_1, out_of_19_2, out_of_19_3, out_of_19_4, out_of_19_5, out_of_19_6, out_of_19_7, out_of_19_8, out_of_19_9, out_of_19_10, out_of_19_11, out_of_19_12, out_of_19_13, out_of_19_14, out_of_19_15, out_of_19_16, out_of_19_17, out_of_19_18, out_of_19_19, out_of_19_20, out_of_19_21, out_of_19_22, out_of_19_23, out_of_19_24, out_of_19_25, out_of_19_26, out_of_19_27, out_of_19_28, out_of_19_29, out_of_19_30, out_of_19_31, out_of_20_0, out_of_20_1, out_of_20_2, out_of_20_3, out_of_20_4, out_of_20_5, out_of_20_6, out_of_20_7, out_of_20_8, out_of_20_9, out_of_20_10, out_of_20_11, out_of_20_12, out_of_20_13, out_of_20_14, out_of_20_15, out_of_20_16, out_of_20_17, out_of_20_18, out_of_20_19, out_of_20_20, out_of_20_21, out_of_20_22, out_of_20_23, out_of_20_24, out_of_20_25, out_of_20_26, out_of_20_27, out_of_20_28, out_of_20_29, out_of_20_30, out_of_20_31, out_of_21_0, out_of_21_1, out_of_21_2, out_of_21_3, out_of_21_4, out_of_21_5, out_of_21_6, out_of_21_7, out_of_21_8, out_of_21_9, out_of_21_10, out_of_21_11, out_of_21_12, out_of_21_13, out_of_21_14, out_of_21_15, out_of_21_16, out_of_21_17, out_of_21_18, out_of_21_19, out_of_21_20, out_of_21_21, out_of_21_22, out_of_21_23, out_of_21_24, out_of_21_25, out_of_21_26, out_of_21_27, out_of_21_28, out_of_21_29, out_of_21_30, out_of_21_31, out_of_22_0, out_of_22_1, out_of_22_2, out_of_22_3, out_of_22_4, out_of_22_5, out_of_22_6, out_of_22_7, out_of_22_8, out_of_22_9, out_of_22_10, out_of_22_11, out_of_22_12, out_of_22_13, out_of_22_14, out_of_22_15, out_of_22_16, out_of_22_17, out_of_22_18, out_of_22_19, out_of_22_20, out_of_22_21, out_of_22_22, out_of_22_23, out_of_22_24, out_of_22_25, out_of_22_26, out_of_22_27, out_of_22_28, out_of_22_29, out_of_22_30, out_of_22_31, out_of_23_0, out_of_23_1, out_of_23_2, out_of_23_3, out_of_23_4, out_of_23_5, out_of_23_6, out_of_23_7, out_of_23_8, out_of_23_9, out_of_23_10, out_of_23_11, out_of_23_12, out_of_23_13, out_of_23_14, out_of_23_15, out_of_23_16, out_of_23_17, out_of_23_18, out_of_23_19, out_of_23_20, out_of_23_21, out_of_23_22, out_of_23_23, out_of_23_24, out_of_23_25, out_of_23_26, out_of_23_27, out_of_23_28, out_of_23_29, out_of_23_30, out_of_23_31, out_of_24_0, out_of_24_1, out_of_24_2, out_of_24_3, out_of_24_4, out_of_24_5, out_of_24_6, out_of_24_7, out_of_24_8, out_of_24_9, out_of_24_10, out_of_24_11, out_of_24_12, out_of_24_13, out_of_24_14, out_of_24_15, out_of_24_16, out_of_24_17, out_of_24_18, out_of_24_19, out_of_24_20, out_of_24_21, out_of_24_22, out_of_24_23, out_of_24_24, out_of_24_25, out_of_24_26, out_of_24_27, out_of_24_28, out_of_24_29, out_of_24_30, out_of_24_31, out_of_25_0, out_of_25_1, out_of_25_2, out_of_25_3, out_of_25_4, out_of_25_5, out_of_25_6, out_of_25_7, out_of_25_8, out_of_25_9, out_of_25_10, out_of_25_11, out_of_25_12, out_of_25_13, out_of_25_14, out_of_25_15, out_of_25_16, out_of_25_17, out_of_25_18, out_of_25_19, out_of_25_20, out_of_25_21, out_of_25_22, out_of_25_23, out_of_25_24, out_of_25_25, out_of_25_26, out_of_25_27, out_of_25_28, out_of_25_29, out_of_25_30, out_of_25_31, out_of_26_0, out_of_26_1, out_of_26_2, out_of_26_3, out_of_26_4, out_of_26_5, out_of_26_6, out_of_26_7, out_of_26_8, out_of_26_9, out_of_26_10, out_of_26_11, out_of_26_12, out_of_26_13, out_of_26_14, out_of_26_15, out_of_26_16, out_of_26_17, out_of_26_18, out_of_26_19, out_of_26_20, out_of_26_21, out_of_26_22, out_of_26_23, out_of_26_24, out_of_26_25, out_of_26_26, out_of_26_27, out_of_26_28, out_of_26_29, out_of_26_30, out_of_26_31, out_of_27_0, out_of_27_1, out_of_27_2, out_of_27_3, out_of_27_4, out_of_27_5, out_of_27_6, out_of_27_7, out_of_27_8, out_of_27_9, out_of_27_10, out_of_27_11, out_of_27_12, out_of_27_13, out_of_27_14, out_of_27_15, out_of_27_16, out_of_27_17, out_of_27_18, out_of_27_19, out_of_27_20, out_of_27_21, out_of_27_22, out_of_27_23, out_of_27_24, out_of_27_25, out_of_27_26, out_of_27_27, out_of_27_28, out_of_27_29, out_of_27_30, out_of_27_31, out_of_28_0, out_of_28_1, out_of_28_2, out_of_28_3, out_of_28_4, out_of_28_5, out_of_28_6, out_of_28_7, out_of_28_8, out_of_28_9, out_of_28_10, out_of_28_11, out_of_28_12, out_of_28_13, out_of_28_14, out_of_28_15, out_of_28_16, out_of_28_17, out_of_28_18, out_of_28_19, out_of_28_20, out_of_28_21, out_of_28_22, out_of_28_23, out_of_28_24, out_of_28_25, out_of_28_26, out_of_28_27, out_of_28_28, out_of_28_29, out_of_28_30, out_of_28_31, out_of_29_0, out_of_29_1, out_of_29_2, out_of_29_3, out_of_29_4, out_of_29_5, out_of_29_6, out_of_29_7, out_of_29_8, out_of_29_9, out_of_29_10, out_of_29_11, out_of_29_12, out_of_29_13, out_of_29_14, out_of_29_15, out_of_29_16, out_of_29_17, out_of_29_18, out_of_29_19, out_of_29_20, out_of_29_21, out_of_29_22, out_of_29_23, out_of_29_24, out_of_29_25, out_of_29_26, out_of_29_27, out_of_29_28, out_of_29_29, out_of_29_30, out_of_29_31, out_of_30_0, out_of_30_1, out_of_30_2, out_of_30_3, out_of_30_4, out_of_30_5, out_of_30_6, out_of_30_7, out_of_30_8, out_of_30_9, out_of_30_10, out_of_30_11, out_of_30_12, out_of_30_13, out_of_30_14, out_of_30_15, out_of_30_16, out_of_30_17, out_of_30_18, out_of_30_19, out_of_30_20, out_of_30_21, out_of_30_22, out_of_30_23, out_of_30_24, out_of_30_25, out_of_30_26, out_of_30_27, out_of_30_28, out_of_30_29, out_of_30_30, out_of_30_31, out_of_31_0, out_of_31_1, out_of_31_2, out_of_31_3, out_of_31_4, out_of_31_5, out_of_31_6, out_of_31_7, out_of_31_8, out_of_31_9, out_of_31_10, out_of_31_11, out_of_31_12, out_of_31_13, out_of_31_14, out_of_31_15, out_of_31_16, out_of_31_17, out_of_31_18, out_of_31_19, out_of_31_20, out_of_31_21, out_of_31_22, out_of_31_23, out_of_31_24, out_of_31_25, out_of_31_26, out_of_31_27, out_of_31_28, out_of_31_29, out_of_31_30, out_of_31_31;

assign {in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27, in_28, in_29, in_30, in_31} = in_buffer;

transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_0(clock, reset, enable, direction, in_31, in_0, out_of_0_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_1(clock, reset, enable, direction, in_30, out_of_0_0, out_of_0_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_2(clock, reset, enable, direction, in_29, out_of_0_1, out_of_0_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_3(clock, reset, enable, direction, in_28, out_of_0_2, out_of_0_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_4(clock, reset, enable, direction, in_27, out_of_0_3, out_of_0_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_5(clock, reset, enable, direction, in_26, out_of_0_4, out_of_0_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_6(clock, reset, enable, direction, in_25, out_of_0_5, out_of_0_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_7(clock, reset, enable, direction, in_24, out_of_0_6, out_of_0_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_8(clock, reset, enable, direction, in_23, out_of_0_7, out_of_0_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_9(clock, reset, enable, direction, in_22, out_of_0_8, out_of_0_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_10(clock, reset, enable, direction, in_21, out_of_0_9, out_of_0_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_11(clock, reset, enable, direction, in_20, out_of_0_10, out_of_0_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_12(clock, reset, enable, direction, in_19, out_of_0_11, out_of_0_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_13(clock, reset, enable, direction, in_18, out_of_0_12, out_of_0_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_14(clock, reset, enable, direction, in_17, out_of_0_13, out_of_0_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_15(clock, reset, enable, direction, in_16, out_of_0_14, out_of_0_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_16(clock, reset, enable, direction, in_15, out_of_0_15, out_of_0_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_17(clock, reset, enable, direction, in_14, out_of_0_16, out_of_0_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_18(clock, reset, enable, direction, in_13, out_of_0_17, out_of_0_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_19(clock, reset, enable, direction, in_12, out_of_0_18, out_of_0_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_20(clock, reset, enable, direction, in_11, out_of_0_19, out_of_0_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_21(clock, reset, enable, direction, in_10, out_of_0_20, out_of_0_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_22(clock, reset, enable, direction, in_9, out_of_0_21, out_of_0_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_23(clock, reset, enable, direction, in_8, out_of_0_22, out_of_0_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_24(clock, reset, enable, direction, in_7, out_of_0_23, out_of_0_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_25(clock, reset, enable, direction, in_6, out_of_0_24, out_of_0_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_26(clock, reset, enable, direction, in_5, out_of_0_25, out_of_0_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_27(clock, reset, enable, direction, in_4, out_of_0_26, out_of_0_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_28(clock, reset, enable, direction, in_3, out_of_0_27, out_of_0_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_29(clock, reset, enable, direction, in_2, out_of_0_28, out_of_0_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_30(clock, reset, enable, direction, in_1, out_of_0_29, out_of_0_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_0_31(clock, reset, enable, direction, in_0, out_of_0_30, out_of_0_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_0(clock, reset, enable, direction, out_of_0_0, in_1, out_of_1_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_1(clock, reset, enable, direction, out_of_0_1, out_of_1_0, out_of_1_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_2(clock, reset, enable, direction, out_of_0_2, out_of_1_1, out_of_1_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_3(clock, reset, enable, direction, out_of_0_3, out_of_1_2, out_of_1_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_4(clock, reset, enable, direction, out_of_0_4, out_of_1_3, out_of_1_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_5(clock, reset, enable, direction, out_of_0_5, out_of_1_4, out_of_1_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_6(clock, reset, enable, direction, out_of_0_6, out_of_1_5, out_of_1_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_7(clock, reset, enable, direction, out_of_0_7, out_of_1_6, out_of_1_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_8(clock, reset, enable, direction, out_of_0_8, out_of_1_7, out_of_1_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_9(clock, reset, enable, direction, out_of_0_9, out_of_1_8, out_of_1_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_10(clock, reset, enable, direction, out_of_0_10, out_of_1_9, out_of_1_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_11(clock, reset, enable, direction, out_of_0_11, out_of_1_10, out_of_1_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_12(clock, reset, enable, direction, out_of_0_12, out_of_1_11, out_of_1_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_13(clock, reset, enable, direction, out_of_0_13, out_of_1_12, out_of_1_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_14(clock, reset, enable, direction, out_of_0_14, out_of_1_13, out_of_1_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_15(clock, reset, enable, direction, out_of_0_15, out_of_1_14, out_of_1_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_16(clock, reset, enable, direction, out_of_0_16, out_of_1_15, out_of_1_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_17(clock, reset, enable, direction, out_of_0_17, out_of_1_16, out_of_1_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_18(clock, reset, enable, direction, out_of_0_18, out_of_1_17, out_of_1_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_19(clock, reset, enable, direction, out_of_0_19, out_of_1_18, out_of_1_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_20(clock, reset, enable, direction, out_of_0_20, out_of_1_19, out_of_1_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_21(clock, reset, enable, direction, out_of_0_21, out_of_1_20, out_of_1_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_22(clock, reset, enable, direction, out_of_0_22, out_of_1_21, out_of_1_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_23(clock, reset, enable, direction, out_of_0_23, out_of_1_22, out_of_1_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_24(clock, reset, enable, direction, out_of_0_24, out_of_1_23, out_of_1_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_25(clock, reset, enable, direction, out_of_0_25, out_of_1_24, out_of_1_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_26(clock, reset, enable, direction, out_of_0_26, out_of_1_25, out_of_1_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_27(clock, reset, enable, direction, out_of_0_27, out_of_1_26, out_of_1_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_28(clock, reset, enable, direction, out_of_0_28, out_of_1_27, out_of_1_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_29(clock, reset, enable, direction, out_of_0_29, out_of_1_28, out_of_1_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_30(clock, reset, enable, direction, out_of_0_30, out_of_1_29, out_of_1_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_1_31(clock, reset, enable, direction, out_of_0_31, out_of_1_30, out_of_1_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_0(clock, reset, enable, direction, out_of_1_0, in_2, out_of_2_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_1(clock, reset, enable, direction, out_of_1_1, out_of_2_0, out_of_2_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_2(clock, reset, enable, direction, out_of_1_2, out_of_2_1, out_of_2_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_3(clock, reset, enable, direction, out_of_1_3, out_of_2_2, out_of_2_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_4(clock, reset, enable, direction, out_of_1_4, out_of_2_3, out_of_2_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_5(clock, reset, enable, direction, out_of_1_5, out_of_2_4, out_of_2_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_6(clock, reset, enable, direction, out_of_1_6, out_of_2_5, out_of_2_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_7(clock, reset, enable, direction, out_of_1_7, out_of_2_6, out_of_2_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_8(clock, reset, enable, direction, out_of_1_8, out_of_2_7, out_of_2_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_9(clock, reset, enable, direction, out_of_1_9, out_of_2_8, out_of_2_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_10(clock, reset, enable, direction, out_of_1_10, out_of_2_9, out_of_2_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_11(clock, reset, enable, direction, out_of_1_11, out_of_2_10, out_of_2_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_12(clock, reset, enable, direction, out_of_1_12, out_of_2_11, out_of_2_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_13(clock, reset, enable, direction, out_of_1_13, out_of_2_12, out_of_2_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_14(clock, reset, enable, direction, out_of_1_14, out_of_2_13, out_of_2_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_15(clock, reset, enable, direction, out_of_1_15, out_of_2_14, out_of_2_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_16(clock, reset, enable, direction, out_of_1_16, out_of_2_15, out_of_2_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_17(clock, reset, enable, direction, out_of_1_17, out_of_2_16, out_of_2_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_18(clock, reset, enable, direction, out_of_1_18, out_of_2_17, out_of_2_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_19(clock, reset, enable, direction, out_of_1_19, out_of_2_18, out_of_2_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_20(clock, reset, enable, direction, out_of_1_20, out_of_2_19, out_of_2_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_21(clock, reset, enable, direction, out_of_1_21, out_of_2_20, out_of_2_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_22(clock, reset, enable, direction, out_of_1_22, out_of_2_21, out_of_2_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_23(clock, reset, enable, direction, out_of_1_23, out_of_2_22, out_of_2_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_24(clock, reset, enable, direction, out_of_1_24, out_of_2_23, out_of_2_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_25(clock, reset, enable, direction, out_of_1_25, out_of_2_24, out_of_2_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_26(clock, reset, enable, direction, out_of_1_26, out_of_2_25, out_of_2_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_27(clock, reset, enable, direction, out_of_1_27, out_of_2_26, out_of_2_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_28(clock, reset, enable, direction, out_of_1_28, out_of_2_27, out_of_2_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_29(clock, reset, enable, direction, out_of_1_29, out_of_2_28, out_of_2_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_30(clock, reset, enable, direction, out_of_1_30, out_of_2_29, out_of_2_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_2_31(clock, reset, enable, direction, out_of_1_31, out_of_2_30, out_of_2_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_0(clock, reset, enable, direction, out_of_2_0, in_3, out_of_3_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_1(clock, reset, enable, direction, out_of_2_1, out_of_3_0, out_of_3_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_2(clock, reset, enable, direction, out_of_2_2, out_of_3_1, out_of_3_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_3(clock, reset, enable, direction, out_of_2_3, out_of_3_2, out_of_3_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_4(clock, reset, enable, direction, out_of_2_4, out_of_3_3, out_of_3_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_5(clock, reset, enable, direction, out_of_2_5, out_of_3_4, out_of_3_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_6(clock, reset, enable, direction, out_of_2_6, out_of_3_5, out_of_3_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_7(clock, reset, enable, direction, out_of_2_7, out_of_3_6, out_of_3_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_8(clock, reset, enable, direction, out_of_2_8, out_of_3_7, out_of_3_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_9(clock, reset, enable, direction, out_of_2_9, out_of_3_8, out_of_3_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_10(clock, reset, enable, direction, out_of_2_10, out_of_3_9, out_of_3_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_11(clock, reset, enable, direction, out_of_2_11, out_of_3_10, out_of_3_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_12(clock, reset, enable, direction, out_of_2_12, out_of_3_11, out_of_3_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_13(clock, reset, enable, direction, out_of_2_13, out_of_3_12, out_of_3_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_14(clock, reset, enable, direction, out_of_2_14, out_of_3_13, out_of_3_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_15(clock, reset, enable, direction, out_of_2_15, out_of_3_14, out_of_3_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_16(clock, reset, enable, direction, out_of_2_16, out_of_3_15, out_of_3_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_17(clock, reset, enable, direction, out_of_2_17, out_of_3_16, out_of_3_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_18(clock, reset, enable, direction, out_of_2_18, out_of_3_17, out_of_3_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_19(clock, reset, enable, direction, out_of_2_19, out_of_3_18, out_of_3_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_20(clock, reset, enable, direction, out_of_2_20, out_of_3_19, out_of_3_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_21(clock, reset, enable, direction, out_of_2_21, out_of_3_20, out_of_3_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_22(clock, reset, enable, direction, out_of_2_22, out_of_3_21, out_of_3_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_23(clock, reset, enable, direction, out_of_2_23, out_of_3_22, out_of_3_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_24(clock, reset, enable, direction, out_of_2_24, out_of_3_23, out_of_3_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_25(clock, reset, enable, direction, out_of_2_25, out_of_3_24, out_of_3_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_26(clock, reset, enable, direction, out_of_2_26, out_of_3_25, out_of_3_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_27(clock, reset, enable, direction, out_of_2_27, out_of_3_26, out_of_3_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_28(clock, reset, enable, direction, out_of_2_28, out_of_3_27, out_of_3_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_29(clock, reset, enable, direction, out_of_2_29, out_of_3_28, out_of_3_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_30(clock, reset, enable, direction, out_of_2_30, out_of_3_29, out_of_3_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_3_31(clock, reset, enable, direction, out_of_2_31, out_of_3_30, out_of_3_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_0(clock, reset, enable, direction, out_of_3_0, in_4, out_of_4_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_1(clock, reset, enable, direction, out_of_3_1, out_of_4_0, out_of_4_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_2(clock, reset, enable, direction, out_of_3_2, out_of_4_1, out_of_4_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_3(clock, reset, enable, direction, out_of_3_3, out_of_4_2, out_of_4_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_4(clock, reset, enable, direction, out_of_3_4, out_of_4_3, out_of_4_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_5(clock, reset, enable, direction, out_of_3_5, out_of_4_4, out_of_4_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_6(clock, reset, enable, direction, out_of_3_6, out_of_4_5, out_of_4_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_7(clock, reset, enable, direction, out_of_3_7, out_of_4_6, out_of_4_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_8(clock, reset, enable, direction, out_of_3_8, out_of_4_7, out_of_4_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_9(clock, reset, enable, direction, out_of_3_9, out_of_4_8, out_of_4_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_10(clock, reset, enable, direction, out_of_3_10, out_of_4_9, out_of_4_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_11(clock, reset, enable, direction, out_of_3_11, out_of_4_10, out_of_4_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_12(clock, reset, enable, direction, out_of_3_12, out_of_4_11, out_of_4_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_13(clock, reset, enable, direction, out_of_3_13, out_of_4_12, out_of_4_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_14(clock, reset, enable, direction, out_of_3_14, out_of_4_13, out_of_4_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_15(clock, reset, enable, direction, out_of_3_15, out_of_4_14, out_of_4_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_16(clock, reset, enable, direction, out_of_3_16, out_of_4_15, out_of_4_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_17(clock, reset, enable, direction, out_of_3_17, out_of_4_16, out_of_4_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_18(clock, reset, enable, direction, out_of_3_18, out_of_4_17, out_of_4_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_19(clock, reset, enable, direction, out_of_3_19, out_of_4_18, out_of_4_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_20(clock, reset, enable, direction, out_of_3_20, out_of_4_19, out_of_4_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_21(clock, reset, enable, direction, out_of_3_21, out_of_4_20, out_of_4_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_22(clock, reset, enable, direction, out_of_3_22, out_of_4_21, out_of_4_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_23(clock, reset, enable, direction, out_of_3_23, out_of_4_22, out_of_4_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_24(clock, reset, enable, direction, out_of_3_24, out_of_4_23, out_of_4_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_25(clock, reset, enable, direction, out_of_3_25, out_of_4_24, out_of_4_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_26(clock, reset, enable, direction, out_of_3_26, out_of_4_25, out_of_4_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_27(clock, reset, enable, direction, out_of_3_27, out_of_4_26, out_of_4_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_28(clock, reset, enable, direction, out_of_3_28, out_of_4_27, out_of_4_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_29(clock, reset, enable, direction, out_of_3_29, out_of_4_28, out_of_4_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_30(clock, reset, enable, direction, out_of_3_30, out_of_4_29, out_of_4_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_4_31(clock, reset, enable, direction, out_of_3_31, out_of_4_30, out_of_4_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_0(clock, reset, enable, direction, out_of_4_0, in_5, out_of_5_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_1(clock, reset, enable, direction, out_of_4_1, out_of_5_0, out_of_5_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_2(clock, reset, enable, direction, out_of_4_2, out_of_5_1, out_of_5_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_3(clock, reset, enable, direction, out_of_4_3, out_of_5_2, out_of_5_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_4(clock, reset, enable, direction, out_of_4_4, out_of_5_3, out_of_5_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_5(clock, reset, enable, direction, out_of_4_5, out_of_5_4, out_of_5_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_6(clock, reset, enable, direction, out_of_4_6, out_of_5_5, out_of_5_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_7(clock, reset, enable, direction, out_of_4_7, out_of_5_6, out_of_5_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_8(clock, reset, enable, direction, out_of_4_8, out_of_5_7, out_of_5_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_9(clock, reset, enable, direction, out_of_4_9, out_of_5_8, out_of_5_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_10(clock, reset, enable, direction, out_of_4_10, out_of_5_9, out_of_5_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_11(clock, reset, enable, direction, out_of_4_11, out_of_5_10, out_of_5_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_12(clock, reset, enable, direction, out_of_4_12, out_of_5_11, out_of_5_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_13(clock, reset, enable, direction, out_of_4_13, out_of_5_12, out_of_5_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_14(clock, reset, enable, direction, out_of_4_14, out_of_5_13, out_of_5_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_15(clock, reset, enable, direction, out_of_4_15, out_of_5_14, out_of_5_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_16(clock, reset, enable, direction, out_of_4_16, out_of_5_15, out_of_5_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_17(clock, reset, enable, direction, out_of_4_17, out_of_5_16, out_of_5_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_18(clock, reset, enable, direction, out_of_4_18, out_of_5_17, out_of_5_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_19(clock, reset, enable, direction, out_of_4_19, out_of_5_18, out_of_5_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_20(clock, reset, enable, direction, out_of_4_20, out_of_5_19, out_of_5_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_21(clock, reset, enable, direction, out_of_4_21, out_of_5_20, out_of_5_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_22(clock, reset, enable, direction, out_of_4_22, out_of_5_21, out_of_5_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_23(clock, reset, enable, direction, out_of_4_23, out_of_5_22, out_of_5_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_24(clock, reset, enable, direction, out_of_4_24, out_of_5_23, out_of_5_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_25(clock, reset, enable, direction, out_of_4_25, out_of_5_24, out_of_5_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_26(clock, reset, enable, direction, out_of_4_26, out_of_5_25, out_of_5_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_27(clock, reset, enable, direction, out_of_4_27, out_of_5_26, out_of_5_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_28(clock, reset, enable, direction, out_of_4_28, out_of_5_27, out_of_5_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_29(clock, reset, enable, direction, out_of_4_29, out_of_5_28, out_of_5_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_30(clock, reset, enable, direction, out_of_4_30, out_of_5_29, out_of_5_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_5_31(clock, reset, enable, direction, out_of_4_31, out_of_5_30, out_of_5_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_0(clock, reset, enable, direction, out_of_5_0, in_6, out_of_6_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_1(clock, reset, enable, direction, out_of_5_1, out_of_6_0, out_of_6_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_2(clock, reset, enable, direction, out_of_5_2, out_of_6_1, out_of_6_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_3(clock, reset, enable, direction, out_of_5_3, out_of_6_2, out_of_6_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_4(clock, reset, enable, direction, out_of_5_4, out_of_6_3, out_of_6_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_5(clock, reset, enable, direction, out_of_5_5, out_of_6_4, out_of_6_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_6(clock, reset, enable, direction, out_of_5_6, out_of_6_5, out_of_6_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_7(clock, reset, enable, direction, out_of_5_7, out_of_6_6, out_of_6_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_8(clock, reset, enable, direction, out_of_5_8, out_of_6_7, out_of_6_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_9(clock, reset, enable, direction, out_of_5_9, out_of_6_8, out_of_6_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_10(clock, reset, enable, direction, out_of_5_10, out_of_6_9, out_of_6_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_11(clock, reset, enable, direction, out_of_5_11, out_of_6_10, out_of_6_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_12(clock, reset, enable, direction, out_of_5_12, out_of_6_11, out_of_6_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_13(clock, reset, enable, direction, out_of_5_13, out_of_6_12, out_of_6_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_14(clock, reset, enable, direction, out_of_5_14, out_of_6_13, out_of_6_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_15(clock, reset, enable, direction, out_of_5_15, out_of_6_14, out_of_6_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_16(clock, reset, enable, direction, out_of_5_16, out_of_6_15, out_of_6_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_17(clock, reset, enable, direction, out_of_5_17, out_of_6_16, out_of_6_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_18(clock, reset, enable, direction, out_of_5_18, out_of_6_17, out_of_6_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_19(clock, reset, enable, direction, out_of_5_19, out_of_6_18, out_of_6_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_20(clock, reset, enable, direction, out_of_5_20, out_of_6_19, out_of_6_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_21(clock, reset, enable, direction, out_of_5_21, out_of_6_20, out_of_6_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_22(clock, reset, enable, direction, out_of_5_22, out_of_6_21, out_of_6_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_23(clock, reset, enable, direction, out_of_5_23, out_of_6_22, out_of_6_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_24(clock, reset, enable, direction, out_of_5_24, out_of_6_23, out_of_6_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_25(clock, reset, enable, direction, out_of_5_25, out_of_6_24, out_of_6_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_26(clock, reset, enable, direction, out_of_5_26, out_of_6_25, out_of_6_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_27(clock, reset, enable, direction, out_of_5_27, out_of_6_26, out_of_6_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_28(clock, reset, enable, direction, out_of_5_28, out_of_6_27, out_of_6_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_29(clock, reset, enable, direction, out_of_5_29, out_of_6_28, out_of_6_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_30(clock, reset, enable, direction, out_of_5_30, out_of_6_29, out_of_6_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_6_31(clock, reset, enable, direction, out_of_5_31, out_of_6_30, out_of_6_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_0(clock, reset, enable, direction, out_of_6_0, in_7, out_of_7_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_1(clock, reset, enable, direction, out_of_6_1, out_of_7_0, out_of_7_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_2(clock, reset, enable, direction, out_of_6_2, out_of_7_1, out_of_7_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_3(clock, reset, enable, direction, out_of_6_3, out_of_7_2, out_of_7_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_4(clock, reset, enable, direction, out_of_6_4, out_of_7_3, out_of_7_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_5(clock, reset, enable, direction, out_of_6_5, out_of_7_4, out_of_7_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_6(clock, reset, enable, direction, out_of_6_6, out_of_7_5, out_of_7_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_7(clock, reset, enable, direction, out_of_6_7, out_of_7_6, out_of_7_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_8(clock, reset, enable, direction, out_of_6_8, out_of_7_7, out_of_7_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_9(clock, reset, enable, direction, out_of_6_9, out_of_7_8, out_of_7_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_10(clock, reset, enable, direction, out_of_6_10, out_of_7_9, out_of_7_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_11(clock, reset, enable, direction, out_of_6_11, out_of_7_10, out_of_7_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_12(clock, reset, enable, direction, out_of_6_12, out_of_7_11, out_of_7_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_13(clock, reset, enable, direction, out_of_6_13, out_of_7_12, out_of_7_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_14(clock, reset, enable, direction, out_of_6_14, out_of_7_13, out_of_7_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_15(clock, reset, enable, direction, out_of_6_15, out_of_7_14, out_of_7_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_16(clock, reset, enable, direction, out_of_6_16, out_of_7_15, out_of_7_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_17(clock, reset, enable, direction, out_of_6_17, out_of_7_16, out_of_7_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_18(clock, reset, enable, direction, out_of_6_18, out_of_7_17, out_of_7_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_19(clock, reset, enable, direction, out_of_6_19, out_of_7_18, out_of_7_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_20(clock, reset, enable, direction, out_of_6_20, out_of_7_19, out_of_7_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_21(clock, reset, enable, direction, out_of_6_21, out_of_7_20, out_of_7_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_22(clock, reset, enable, direction, out_of_6_22, out_of_7_21, out_of_7_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_23(clock, reset, enable, direction, out_of_6_23, out_of_7_22, out_of_7_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_24(clock, reset, enable, direction, out_of_6_24, out_of_7_23, out_of_7_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_25(clock, reset, enable, direction, out_of_6_25, out_of_7_24, out_of_7_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_26(clock, reset, enable, direction, out_of_6_26, out_of_7_25, out_of_7_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_27(clock, reset, enable, direction, out_of_6_27, out_of_7_26, out_of_7_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_28(clock, reset, enable, direction, out_of_6_28, out_of_7_27, out_of_7_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_29(clock, reset, enable, direction, out_of_6_29, out_of_7_28, out_of_7_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_30(clock, reset, enable, direction, out_of_6_30, out_of_7_29, out_of_7_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_7_31(clock, reset, enable, direction, out_of_6_31, out_of_7_30, out_of_7_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_0(clock, reset, enable, direction, out_of_7_0, in_8, out_of_8_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_1(clock, reset, enable, direction, out_of_7_1, out_of_8_0, out_of_8_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_2(clock, reset, enable, direction, out_of_7_2, out_of_8_1, out_of_8_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_3(clock, reset, enable, direction, out_of_7_3, out_of_8_2, out_of_8_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_4(clock, reset, enable, direction, out_of_7_4, out_of_8_3, out_of_8_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_5(clock, reset, enable, direction, out_of_7_5, out_of_8_4, out_of_8_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_6(clock, reset, enable, direction, out_of_7_6, out_of_8_5, out_of_8_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_7(clock, reset, enable, direction, out_of_7_7, out_of_8_6, out_of_8_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_8(clock, reset, enable, direction, out_of_7_8, out_of_8_7, out_of_8_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_9(clock, reset, enable, direction, out_of_7_9, out_of_8_8, out_of_8_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_10(clock, reset, enable, direction, out_of_7_10, out_of_8_9, out_of_8_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_11(clock, reset, enable, direction, out_of_7_11, out_of_8_10, out_of_8_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_12(clock, reset, enable, direction, out_of_7_12, out_of_8_11, out_of_8_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_13(clock, reset, enable, direction, out_of_7_13, out_of_8_12, out_of_8_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_14(clock, reset, enable, direction, out_of_7_14, out_of_8_13, out_of_8_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_15(clock, reset, enable, direction, out_of_7_15, out_of_8_14, out_of_8_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_16(clock, reset, enable, direction, out_of_7_16, out_of_8_15, out_of_8_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_17(clock, reset, enable, direction, out_of_7_17, out_of_8_16, out_of_8_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_18(clock, reset, enable, direction, out_of_7_18, out_of_8_17, out_of_8_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_19(clock, reset, enable, direction, out_of_7_19, out_of_8_18, out_of_8_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_20(clock, reset, enable, direction, out_of_7_20, out_of_8_19, out_of_8_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_21(clock, reset, enable, direction, out_of_7_21, out_of_8_20, out_of_8_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_22(clock, reset, enable, direction, out_of_7_22, out_of_8_21, out_of_8_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_23(clock, reset, enable, direction, out_of_7_23, out_of_8_22, out_of_8_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_24(clock, reset, enable, direction, out_of_7_24, out_of_8_23, out_of_8_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_25(clock, reset, enable, direction, out_of_7_25, out_of_8_24, out_of_8_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_26(clock, reset, enable, direction, out_of_7_26, out_of_8_25, out_of_8_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_27(clock, reset, enable, direction, out_of_7_27, out_of_8_26, out_of_8_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_28(clock, reset, enable, direction, out_of_7_28, out_of_8_27, out_of_8_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_29(clock, reset, enable, direction, out_of_7_29, out_of_8_28, out_of_8_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_30(clock, reset, enable, direction, out_of_7_30, out_of_8_29, out_of_8_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_8_31(clock, reset, enable, direction, out_of_7_31, out_of_8_30, out_of_8_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_0(clock, reset, enable, direction, out_of_8_0, in_9, out_of_9_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_1(clock, reset, enable, direction, out_of_8_1, out_of_9_0, out_of_9_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_2(clock, reset, enable, direction, out_of_8_2, out_of_9_1, out_of_9_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_3(clock, reset, enable, direction, out_of_8_3, out_of_9_2, out_of_9_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_4(clock, reset, enable, direction, out_of_8_4, out_of_9_3, out_of_9_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_5(clock, reset, enable, direction, out_of_8_5, out_of_9_4, out_of_9_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_6(clock, reset, enable, direction, out_of_8_6, out_of_9_5, out_of_9_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_7(clock, reset, enable, direction, out_of_8_7, out_of_9_6, out_of_9_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_8(clock, reset, enable, direction, out_of_8_8, out_of_9_7, out_of_9_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_9(clock, reset, enable, direction, out_of_8_9, out_of_9_8, out_of_9_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_10(clock, reset, enable, direction, out_of_8_10, out_of_9_9, out_of_9_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_11(clock, reset, enable, direction, out_of_8_11, out_of_9_10, out_of_9_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_12(clock, reset, enable, direction, out_of_8_12, out_of_9_11, out_of_9_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_13(clock, reset, enable, direction, out_of_8_13, out_of_9_12, out_of_9_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_14(clock, reset, enable, direction, out_of_8_14, out_of_9_13, out_of_9_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_15(clock, reset, enable, direction, out_of_8_15, out_of_9_14, out_of_9_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_16(clock, reset, enable, direction, out_of_8_16, out_of_9_15, out_of_9_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_17(clock, reset, enable, direction, out_of_8_17, out_of_9_16, out_of_9_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_18(clock, reset, enable, direction, out_of_8_18, out_of_9_17, out_of_9_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_19(clock, reset, enable, direction, out_of_8_19, out_of_9_18, out_of_9_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_20(clock, reset, enable, direction, out_of_8_20, out_of_9_19, out_of_9_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_21(clock, reset, enable, direction, out_of_8_21, out_of_9_20, out_of_9_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_22(clock, reset, enable, direction, out_of_8_22, out_of_9_21, out_of_9_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_23(clock, reset, enable, direction, out_of_8_23, out_of_9_22, out_of_9_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_24(clock, reset, enable, direction, out_of_8_24, out_of_9_23, out_of_9_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_25(clock, reset, enable, direction, out_of_8_25, out_of_9_24, out_of_9_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_26(clock, reset, enable, direction, out_of_8_26, out_of_9_25, out_of_9_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_27(clock, reset, enable, direction, out_of_8_27, out_of_9_26, out_of_9_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_28(clock, reset, enable, direction, out_of_8_28, out_of_9_27, out_of_9_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_29(clock, reset, enable, direction, out_of_8_29, out_of_9_28, out_of_9_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_30(clock, reset, enable, direction, out_of_8_30, out_of_9_29, out_of_9_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_9_31(clock, reset, enable, direction, out_of_8_31, out_of_9_30, out_of_9_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_0(clock, reset, enable, direction, out_of_9_0, in_10, out_of_10_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_1(clock, reset, enable, direction, out_of_9_1, out_of_10_0, out_of_10_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_2(clock, reset, enable, direction, out_of_9_2, out_of_10_1, out_of_10_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_3(clock, reset, enable, direction, out_of_9_3, out_of_10_2, out_of_10_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_4(clock, reset, enable, direction, out_of_9_4, out_of_10_3, out_of_10_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_5(clock, reset, enable, direction, out_of_9_5, out_of_10_4, out_of_10_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_6(clock, reset, enable, direction, out_of_9_6, out_of_10_5, out_of_10_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_7(clock, reset, enable, direction, out_of_9_7, out_of_10_6, out_of_10_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_8(clock, reset, enable, direction, out_of_9_8, out_of_10_7, out_of_10_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_9(clock, reset, enable, direction, out_of_9_9, out_of_10_8, out_of_10_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_10(clock, reset, enable, direction, out_of_9_10, out_of_10_9, out_of_10_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_11(clock, reset, enable, direction, out_of_9_11, out_of_10_10, out_of_10_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_12(clock, reset, enable, direction, out_of_9_12, out_of_10_11, out_of_10_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_13(clock, reset, enable, direction, out_of_9_13, out_of_10_12, out_of_10_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_14(clock, reset, enable, direction, out_of_9_14, out_of_10_13, out_of_10_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_15(clock, reset, enable, direction, out_of_9_15, out_of_10_14, out_of_10_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_16(clock, reset, enable, direction, out_of_9_16, out_of_10_15, out_of_10_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_17(clock, reset, enable, direction, out_of_9_17, out_of_10_16, out_of_10_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_18(clock, reset, enable, direction, out_of_9_18, out_of_10_17, out_of_10_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_19(clock, reset, enable, direction, out_of_9_19, out_of_10_18, out_of_10_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_20(clock, reset, enable, direction, out_of_9_20, out_of_10_19, out_of_10_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_21(clock, reset, enable, direction, out_of_9_21, out_of_10_20, out_of_10_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_22(clock, reset, enable, direction, out_of_9_22, out_of_10_21, out_of_10_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_23(clock, reset, enable, direction, out_of_9_23, out_of_10_22, out_of_10_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_24(clock, reset, enable, direction, out_of_9_24, out_of_10_23, out_of_10_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_25(clock, reset, enable, direction, out_of_9_25, out_of_10_24, out_of_10_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_26(clock, reset, enable, direction, out_of_9_26, out_of_10_25, out_of_10_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_27(clock, reset, enable, direction, out_of_9_27, out_of_10_26, out_of_10_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_28(clock, reset, enable, direction, out_of_9_28, out_of_10_27, out_of_10_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_29(clock, reset, enable, direction, out_of_9_29, out_of_10_28, out_of_10_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_30(clock, reset, enable, direction, out_of_9_30, out_of_10_29, out_of_10_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_10_31(clock, reset, enable, direction, out_of_9_31, out_of_10_30, out_of_10_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_0(clock, reset, enable, direction, out_of_10_0, in_11, out_of_11_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_1(clock, reset, enable, direction, out_of_10_1, out_of_11_0, out_of_11_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_2(clock, reset, enable, direction, out_of_10_2, out_of_11_1, out_of_11_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_3(clock, reset, enable, direction, out_of_10_3, out_of_11_2, out_of_11_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_4(clock, reset, enable, direction, out_of_10_4, out_of_11_3, out_of_11_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_5(clock, reset, enable, direction, out_of_10_5, out_of_11_4, out_of_11_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_6(clock, reset, enable, direction, out_of_10_6, out_of_11_5, out_of_11_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_7(clock, reset, enable, direction, out_of_10_7, out_of_11_6, out_of_11_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_8(clock, reset, enable, direction, out_of_10_8, out_of_11_7, out_of_11_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_9(clock, reset, enable, direction, out_of_10_9, out_of_11_8, out_of_11_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_10(clock, reset, enable, direction, out_of_10_10, out_of_11_9, out_of_11_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_11(clock, reset, enable, direction, out_of_10_11, out_of_11_10, out_of_11_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_12(clock, reset, enable, direction, out_of_10_12, out_of_11_11, out_of_11_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_13(clock, reset, enable, direction, out_of_10_13, out_of_11_12, out_of_11_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_14(clock, reset, enable, direction, out_of_10_14, out_of_11_13, out_of_11_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_15(clock, reset, enable, direction, out_of_10_15, out_of_11_14, out_of_11_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_16(clock, reset, enable, direction, out_of_10_16, out_of_11_15, out_of_11_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_17(clock, reset, enable, direction, out_of_10_17, out_of_11_16, out_of_11_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_18(clock, reset, enable, direction, out_of_10_18, out_of_11_17, out_of_11_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_19(clock, reset, enable, direction, out_of_10_19, out_of_11_18, out_of_11_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_20(clock, reset, enable, direction, out_of_10_20, out_of_11_19, out_of_11_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_21(clock, reset, enable, direction, out_of_10_21, out_of_11_20, out_of_11_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_22(clock, reset, enable, direction, out_of_10_22, out_of_11_21, out_of_11_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_23(clock, reset, enable, direction, out_of_10_23, out_of_11_22, out_of_11_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_24(clock, reset, enable, direction, out_of_10_24, out_of_11_23, out_of_11_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_25(clock, reset, enable, direction, out_of_10_25, out_of_11_24, out_of_11_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_26(clock, reset, enable, direction, out_of_10_26, out_of_11_25, out_of_11_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_27(clock, reset, enable, direction, out_of_10_27, out_of_11_26, out_of_11_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_28(clock, reset, enable, direction, out_of_10_28, out_of_11_27, out_of_11_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_29(clock, reset, enable, direction, out_of_10_29, out_of_11_28, out_of_11_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_30(clock, reset, enable, direction, out_of_10_30, out_of_11_29, out_of_11_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_11_31(clock, reset, enable, direction, out_of_10_31, out_of_11_30, out_of_11_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_0(clock, reset, enable, direction, out_of_11_0, in_12, out_of_12_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_1(clock, reset, enable, direction, out_of_11_1, out_of_12_0, out_of_12_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_2(clock, reset, enable, direction, out_of_11_2, out_of_12_1, out_of_12_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_3(clock, reset, enable, direction, out_of_11_3, out_of_12_2, out_of_12_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_4(clock, reset, enable, direction, out_of_11_4, out_of_12_3, out_of_12_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_5(clock, reset, enable, direction, out_of_11_5, out_of_12_4, out_of_12_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_6(clock, reset, enable, direction, out_of_11_6, out_of_12_5, out_of_12_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_7(clock, reset, enable, direction, out_of_11_7, out_of_12_6, out_of_12_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_8(clock, reset, enable, direction, out_of_11_8, out_of_12_7, out_of_12_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_9(clock, reset, enable, direction, out_of_11_9, out_of_12_8, out_of_12_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_10(clock, reset, enable, direction, out_of_11_10, out_of_12_9, out_of_12_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_11(clock, reset, enable, direction, out_of_11_11, out_of_12_10, out_of_12_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_12(clock, reset, enable, direction, out_of_11_12, out_of_12_11, out_of_12_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_13(clock, reset, enable, direction, out_of_11_13, out_of_12_12, out_of_12_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_14(clock, reset, enable, direction, out_of_11_14, out_of_12_13, out_of_12_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_15(clock, reset, enable, direction, out_of_11_15, out_of_12_14, out_of_12_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_16(clock, reset, enable, direction, out_of_11_16, out_of_12_15, out_of_12_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_17(clock, reset, enable, direction, out_of_11_17, out_of_12_16, out_of_12_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_18(clock, reset, enable, direction, out_of_11_18, out_of_12_17, out_of_12_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_19(clock, reset, enable, direction, out_of_11_19, out_of_12_18, out_of_12_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_20(clock, reset, enable, direction, out_of_11_20, out_of_12_19, out_of_12_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_21(clock, reset, enable, direction, out_of_11_21, out_of_12_20, out_of_12_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_22(clock, reset, enable, direction, out_of_11_22, out_of_12_21, out_of_12_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_23(clock, reset, enable, direction, out_of_11_23, out_of_12_22, out_of_12_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_24(clock, reset, enable, direction, out_of_11_24, out_of_12_23, out_of_12_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_25(clock, reset, enable, direction, out_of_11_25, out_of_12_24, out_of_12_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_26(clock, reset, enable, direction, out_of_11_26, out_of_12_25, out_of_12_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_27(clock, reset, enable, direction, out_of_11_27, out_of_12_26, out_of_12_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_28(clock, reset, enable, direction, out_of_11_28, out_of_12_27, out_of_12_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_29(clock, reset, enable, direction, out_of_11_29, out_of_12_28, out_of_12_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_30(clock, reset, enable, direction, out_of_11_30, out_of_12_29, out_of_12_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_12_31(clock, reset, enable, direction, out_of_11_31, out_of_12_30, out_of_12_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_0(clock, reset, enable, direction, out_of_12_0, in_13, out_of_13_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_1(clock, reset, enable, direction, out_of_12_1, out_of_13_0, out_of_13_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_2(clock, reset, enable, direction, out_of_12_2, out_of_13_1, out_of_13_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_3(clock, reset, enable, direction, out_of_12_3, out_of_13_2, out_of_13_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_4(clock, reset, enable, direction, out_of_12_4, out_of_13_3, out_of_13_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_5(clock, reset, enable, direction, out_of_12_5, out_of_13_4, out_of_13_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_6(clock, reset, enable, direction, out_of_12_6, out_of_13_5, out_of_13_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_7(clock, reset, enable, direction, out_of_12_7, out_of_13_6, out_of_13_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_8(clock, reset, enable, direction, out_of_12_8, out_of_13_7, out_of_13_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_9(clock, reset, enable, direction, out_of_12_9, out_of_13_8, out_of_13_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_10(clock, reset, enable, direction, out_of_12_10, out_of_13_9, out_of_13_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_11(clock, reset, enable, direction, out_of_12_11, out_of_13_10, out_of_13_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_12(clock, reset, enable, direction, out_of_12_12, out_of_13_11, out_of_13_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_13(clock, reset, enable, direction, out_of_12_13, out_of_13_12, out_of_13_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_14(clock, reset, enable, direction, out_of_12_14, out_of_13_13, out_of_13_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_15(clock, reset, enable, direction, out_of_12_15, out_of_13_14, out_of_13_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_16(clock, reset, enable, direction, out_of_12_16, out_of_13_15, out_of_13_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_17(clock, reset, enable, direction, out_of_12_17, out_of_13_16, out_of_13_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_18(clock, reset, enable, direction, out_of_12_18, out_of_13_17, out_of_13_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_19(clock, reset, enable, direction, out_of_12_19, out_of_13_18, out_of_13_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_20(clock, reset, enable, direction, out_of_12_20, out_of_13_19, out_of_13_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_21(clock, reset, enable, direction, out_of_12_21, out_of_13_20, out_of_13_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_22(clock, reset, enable, direction, out_of_12_22, out_of_13_21, out_of_13_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_23(clock, reset, enable, direction, out_of_12_23, out_of_13_22, out_of_13_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_24(clock, reset, enable, direction, out_of_12_24, out_of_13_23, out_of_13_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_25(clock, reset, enable, direction, out_of_12_25, out_of_13_24, out_of_13_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_26(clock, reset, enable, direction, out_of_12_26, out_of_13_25, out_of_13_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_27(clock, reset, enable, direction, out_of_12_27, out_of_13_26, out_of_13_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_28(clock, reset, enable, direction, out_of_12_28, out_of_13_27, out_of_13_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_29(clock, reset, enable, direction, out_of_12_29, out_of_13_28, out_of_13_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_30(clock, reset, enable, direction, out_of_12_30, out_of_13_29, out_of_13_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_13_31(clock, reset, enable, direction, out_of_12_31, out_of_13_30, out_of_13_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_0(clock, reset, enable, direction, out_of_13_0, in_14, out_of_14_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_1(clock, reset, enable, direction, out_of_13_1, out_of_14_0, out_of_14_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_2(clock, reset, enable, direction, out_of_13_2, out_of_14_1, out_of_14_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_3(clock, reset, enable, direction, out_of_13_3, out_of_14_2, out_of_14_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_4(clock, reset, enable, direction, out_of_13_4, out_of_14_3, out_of_14_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_5(clock, reset, enable, direction, out_of_13_5, out_of_14_4, out_of_14_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_6(clock, reset, enable, direction, out_of_13_6, out_of_14_5, out_of_14_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_7(clock, reset, enable, direction, out_of_13_7, out_of_14_6, out_of_14_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_8(clock, reset, enable, direction, out_of_13_8, out_of_14_7, out_of_14_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_9(clock, reset, enable, direction, out_of_13_9, out_of_14_8, out_of_14_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_10(clock, reset, enable, direction, out_of_13_10, out_of_14_9, out_of_14_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_11(clock, reset, enable, direction, out_of_13_11, out_of_14_10, out_of_14_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_12(clock, reset, enable, direction, out_of_13_12, out_of_14_11, out_of_14_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_13(clock, reset, enable, direction, out_of_13_13, out_of_14_12, out_of_14_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_14(clock, reset, enable, direction, out_of_13_14, out_of_14_13, out_of_14_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_15(clock, reset, enable, direction, out_of_13_15, out_of_14_14, out_of_14_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_16(clock, reset, enable, direction, out_of_13_16, out_of_14_15, out_of_14_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_17(clock, reset, enable, direction, out_of_13_17, out_of_14_16, out_of_14_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_18(clock, reset, enable, direction, out_of_13_18, out_of_14_17, out_of_14_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_19(clock, reset, enable, direction, out_of_13_19, out_of_14_18, out_of_14_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_20(clock, reset, enable, direction, out_of_13_20, out_of_14_19, out_of_14_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_21(clock, reset, enable, direction, out_of_13_21, out_of_14_20, out_of_14_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_22(clock, reset, enable, direction, out_of_13_22, out_of_14_21, out_of_14_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_23(clock, reset, enable, direction, out_of_13_23, out_of_14_22, out_of_14_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_24(clock, reset, enable, direction, out_of_13_24, out_of_14_23, out_of_14_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_25(clock, reset, enable, direction, out_of_13_25, out_of_14_24, out_of_14_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_26(clock, reset, enable, direction, out_of_13_26, out_of_14_25, out_of_14_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_27(clock, reset, enable, direction, out_of_13_27, out_of_14_26, out_of_14_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_28(clock, reset, enable, direction, out_of_13_28, out_of_14_27, out_of_14_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_29(clock, reset, enable, direction, out_of_13_29, out_of_14_28, out_of_14_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_30(clock, reset, enable, direction, out_of_13_30, out_of_14_29, out_of_14_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_14_31(clock, reset, enable, direction, out_of_13_31, out_of_14_30, out_of_14_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_0(clock, reset, enable, direction, out_of_14_0, in_15, out_of_15_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_1(clock, reset, enable, direction, out_of_14_1, out_of_15_0, out_of_15_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_2(clock, reset, enable, direction, out_of_14_2, out_of_15_1, out_of_15_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_3(clock, reset, enable, direction, out_of_14_3, out_of_15_2, out_of_15_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_4(clock, reset, enable, direction, out_of_14_4, out_of_15_3, out_of_15_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_5(clock, reset, enable, direction, out_of_14_5, out_of_15_4, out_of_15_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_6(clock, reset, enable, direction, out_of_14_6, out_of_15_5, out_of_15_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_7(clock, reset, enable, direction, out_of_14_7, out_of_15_6, out_of_15_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_8(clock, reset, enable, direction, out_of_14_8, out_of_15_7, out_of_15_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_9(clock, reset, enable, direction, out_of_14_9, out_of_15_8, out_of_15_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_10(clock, reset, enable, direction, out_of_14_10, out_of_15_9, out_of_15_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_11(clock, reset, enable, direction, out_of_14_11, out_of_15_10, out_of_15_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_12(clock, reset, enable, direction, out_of_14_12, out_of_15_11, out_of_15_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_13(clock, reset, enable, direction, out_of_14_13, out_of_15_12, out_of_15_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_14(clock, reset, enable, direction, out_of_14_14, out_of_15_13, out_of_15_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_15(clock, reset, enable, direction, out_of_14_15, out_of_15_14, out_of_15_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_16(clock, reset, enable, direction, out_of_14_16, out_of_15_15, out_of_15_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_17(clock, reset, enable, direction, out_of_14_17, out_of_15_16, out_of_15_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_18(clock, reset, enable, direction, out_of_14_18, out_of_15_17, out_of_15_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_19(clock, reset, enable, direction, out_of_14_19, out_of_15_18, out_of_15_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_20(clock, reset, enable, direction, out_of_14_20, out_of_15_19, out_of_15_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_21(clock, reset, enable, direction, out_of_14_21, out_of_15_20, out_of_15_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_22(clock, reset, enable, direction, out_of_14_22, out_of_15_21, out_of_15_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_23(clock, reset, enable, direction, out_of_14_23, out_of_15_22, out_of_15_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_24(clock, reset, enable, direction, out_of_14_24, out_of_15_23, out_of_15_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_25(clock, reset, enable, direction, out_of_14_25, out_of_15_24, out_of_15_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_26(clock, reset, enable, direction, out_of_14_26, out_of_15_25, out_of_15_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_27(clock, reset, enable, direction, out_of_14_27, out_of_15_26, out_of_15_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_28(clock, reset, enable, direction, out_of_14_28, out_of_15_27, out_of_15_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_29(clock, reset, enable, direction, out_of_14_29, out_of_15_28, out_of_15_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_30(clock, reset, enable, direction, out_of_14_30, out_of_15_29, out_of_15_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_15_31(clock, reset, enable, direction, out_of_14_31, out_of_15_30, out_of_15_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_0(clock, reset, enable, direction, out_of_15_0, in_16, out_of_16_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_1(clock, reset, enable, direction, out_of_15_1, out_of_16_0, out_of_16_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_2(clock, reset, enable, direction, out_of_15_2, out_of_16_1, out_of_16_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_3(clock, reset, enable, direction, out_of_15_3, out_of_16_2, out_of_16_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_4(clock, reset, enable, direction, out_of_15_4, out_of_16_3, out_of_16_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_5(clock, reset, enable, direction, out_of_15_5, out_of_16_4, out_of_16_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_6(clock, reset, enable, direction, out_of_15_6, out_of_16_5, out_of_16_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_7(clock, reset, enable, direction, out_of_15_7, out_of_16_6, out_of_16_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_8(clock, reset, enable, direction, out_of_15_8, out_of_16_7, out_of_16_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_9(clock, reset, enable, direction, out_of_15_9, out_of_16_8, out_of_16_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_10(clock, reset, enable, direction, out_of_15_10, out_of_16_9, out_of_16_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_11(clock, reset, enable, direction, out_of_15_11, out_of_16_10, out_of_16_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_12(clock, reset, enable, direction, out_of_15_12, out_of_16_11, out_of_16_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_13(clock, reset, enable, direction, out_of_15_13, out_of_16_12, out_of_16_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_14(clock, reset, enable, direction, out_of_15_14, out_of_16_13, out_of_16_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_15(clock, reset, enable, direction, out_of_15_15, out_of_16_14, out_of_16_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_16(clock, reset, enable, direction, out_of_15_16, out_of_16_15, out_of_16_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_17(clock, reset, enable, direction, out_of_15_17, out_of_16_16, out_of_16_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_18(clock, reset, enable, direction, out_of_15_18, out_of_16_17, out_of_16_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_19(clock, reset, enable, direction, out_of_15_19, out_of_16_18, out_of_16_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_20(clock, reset, enable, direction, out_of_15_20, out_of_16_19, out_of_16_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_21(clock, reset, enable, direction, out_of_15_21, out_of_16_20, out_of_16_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_22(clock, reset, enable, direction, out_of_15_22, out_of_16_21, out_of_16_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_23(clock, reset, enable, direction, out_of_15_23, out_of_16_22, out_of_16_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_24(clock, reset, enable, direction, out_of_15_24, out_of_16_23, out_of_16_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_25(clock, reset, enable, direction, out_of_15_25, out_of_16_24, out_of_16_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_26(clock, reset, enable, direction, out_of_15_26, out_of_16_25, out_of_16_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_27(clock, reset, enable, direction, out_of_15_27, out_of_16_26, out_of_16_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_28(clock, reset, enable, direction, out_of_15_28, out_of_16_27, out_of_16_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_29(clock, reset, enable, direction, out_of_15_29, out_of_16_28, out_of_16_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_30(clock, reset, enable, direction, out_of_15_30, out_of_16_29, out_of_16_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_16_31(clock, reset, enable, direction, out_of_15_31, out_of_16_30, out_of_16_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_0(clock, reset, enable, direction, out_of_16_0, in_17, out_of_17_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_1(clock, reset, enable, direction, out_of_16_1, out_of_17_0, out_of_17_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_2(clock, reset, enable, direction, out_of_16_2, out_of_17_1, out_of_17_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_3(clock, reset, enable, direction, out_of_16_3, out_of_17_2, out_of_17_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_4(clock, reset, enable, direction, out_of_16_4, out_of_17_3, out_of_17_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_5(clock, reset, enable, direction, out_of_16_5, out_of_17_4, out_of_17_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_6(clock, reset, enable, direction, out_of_16_6, out_of_17_5, out_of_17_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_7(clock, reset, enable, direction, out_of_16_7, out_of_17_6, out_of_17_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_8(clock, reset, enable, direction, out_of_16_8, out_of_17_7, out_of_17_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_9(clock, reset, enable, direction, out_of_16_9, out_of_17_8, out_of_17_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_10(clock, reset, enable, direction, out_of_16_10, out_of_17_9, out_of_17_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_11(clock, reset, enable, direction, out_of_16_11, out_of_17_10, out_of_17_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_12(clock, reset, enable, direction, out_of_16_12, out_of_17_11, out_of_17_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_13(clock, reset, enable, direction, out_of_16_13, out_of_17_12, out_of_17_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_14(clock, reset, enable, direction, out_of_16_14, out_of_17_13, out_of_17_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_15(clock, reset, enable, direction, out_of_16_15, out_of_17_14, out_of_17_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_16(clock, reset, enable, direction, out_of_16_16, out_of_17_15, out_of_17_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_17(clock, reset, enable, direction, out_of_16_17, out_of_17_16, out_of_17_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_18(clock, reset, enable, direction, out_of_16_18, out_of_17_17, out_of_17_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_19(clock, reset, enable, direction, out_of_16_19, out_of_17_18, out_of_17_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_20(clock, reset, enable, direction, out_of_16_20, out_of_17_19, out_of_17_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_21(clock, reset, enable, direction, out_of_16_21, out_of_17_20, out_of_17_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_22(clock, reset, enable, direction, out_of_16_22, out_of_17_21, out_of_17_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_23(clock, reset, enable, direction, out_of_16_23, out_of_17_22, out_of_17_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_24(clock, reset, enable, direction, out_of_16_24, out_of_17_23, out_of_17_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_25(clock, reset, enable, direction, out_of_16_25, out_of_17_24, out_of_17_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_26(clock, reset, enable, direction, out_of_16_26, out_of_17_25, out_of_17_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_27(clock, reset, enable, direction, out_of_16_27, out_of_17_26, out_of_17_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_28(clock, reset, enable, direction, out_of_16_28, out_of_17_27, out_of_17_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_29(clock, reset, enable, direction, out_of_16_29, out_of_17_28, out_of_17_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_30(clock, reset, enable, direction, out_of_16_30, out_of_17_29, out_of_17_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_17_31(clock, reset, enable, direction, out_of_16_31, out_of_17_30, out_of_17_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_0(clock, reset, enable, direction, out_of_17_0, in_18, out_of_18_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_1(clock, reset, enable, direction, out_of_17_1, out_of_18_0, out_of_18_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_2(clock, reset, enable, direction, out_of_17_2, out_of_18_1, out_of_18_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_3(clock, reset, enable, direction, out_of_17_3, out_of_18_2, out_of_18_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_4(clock, reset, enable, direction, out_of_17_4, out_of_18_3, out_of_18_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_5(clock, reset, enable, direction, out_of_17_5, out_of_18_4, out_of_18_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_6(clock, reset, enable, direction, out_of_17_6, out_of_18_5, out_of_18_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_7(clock, reset, enable, direction, out_of_17_7, out_of_18_6, out_of_18_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_8(clock, reset, enable, direction, out_of_17_8, out_of_18_7, out_of_18_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_9(clock, reset, enable, direction, out_of_17_9, out_of_18_8, out_of_18_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_10(clock, reset, enable, direction, out_of_17_10, out_of_18_9, out_of_18_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_11(clock, reset, enable, direction, out_of_17_11, out_of_18_10, out_of_18_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_12(clock, reset, enable, direction, out_of_17_12, out_of_18_11, out_of_18_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_13(clock, reset, enable, direction, out_of_17_13, out_of_18_12, out_of_18_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_14(clock, reset, enable, direction, out_of_17_14, out_of_18_13, out_of_18_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_15(clock, reset, enable, direction, out_of_17_15, out_of_18_14, out_of_18_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_16(clock, reset, enable, direction, out_of_17_16, out_of_18_15, out_of_18_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_17(clock, reset, enable, direction, out_of_17_17, out_of_18_16, out_of_18_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_18(clock, reset, enable, direction, out_of_17_18, out_of_18_17, out_of_18_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_19(clock, reset, enable, direction, out_of_17_19, out_of_18_18, out_of_18_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_20(clock, reset, enable, direction, out_of_17_20, out_of_18_19, out_of_18_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_21(clock, reset, enable, direction, out_of_17_21, out_of_18_20, out_of_18_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_22(clock, reset, enable, direction, out_of_17_22, out_of_18_21, out_of_18_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_23(clock, reset, enable, direction, out_of_17_23, out_of_18_22, out_of_18_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_24(clock, reset, enable, direction, out_of_17_24, out_of_18_23, out_of_18_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_25(clock, reset, enable, direction, out_of_17_25, out_of_18_24, out_of_18_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_26(clock, reset, enable, direction, out_of_17_26, out_of_18_25, out_of_18_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_27(clock, reset, enable, direction, out_of_17_27, out_of_18_26, out_of_18_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_28(clock, reset, enable, direction, out_of_17_28, out_of_18_27, out_of_18_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_29(clock, reset, enable, direction, out_of_17_29, out_of_18_28, out_of_18_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_30(clock, reset, enable, direction, out_of_17_30, out_of_18_29, out_of_18_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_18_31(clock, reset, enable, direction, out_of_17_31, out_of_18_30, out_of_18_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_0(clock, reset, enable, direction, out_of_18_0, in_19, out_of_19_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_1(clock, reset, enable, direction, out_of_18_1, out_of_19_0, out_of_19_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_2(clock, reset, enable, direction, out_of_18_2, out_of_19_1, out_of_19_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_3(clock, reset, enable, direction, out_of_18_3, out_of_19_2, out_of_19_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_4(clock, reset, enable, direction, out_of_18_4, out_of_19_3, out_of_19_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_5(clock, reset, enable, direction, out_of_18_5, out_of_19_4, out_of_19_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_6(clock, reset, enable, direction, out_of_18_6, out_of_19_5, out_of_19_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_7(clock, reset, enable, direction, out_of_18_7, out_of_19_6, out_of_19_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_8(clock, reset, enable, direction, out_of_18_8, out_of_19_7, out_of_19_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_9(clock, reset, enable, direction, out_of_18_9, out_of_19_8, out_of_19_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_10(clock, reset, enable, direction, out_of_18_10, out_of_19_9, out_of_19_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_11(clock, reset, enable, direction, out_of_18_11, out_of_19_10, out_of_19_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_12(clock, reset, enable, direction, out_of_18_12, out_of_19_11, out_of_19_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_13(clock, reset, enable, direction, out_of_18_13, out_of_19_12, out_of_19_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_14(clock, reset, enable, direction, out_of_18_14, out_of_19_13, out_of_19_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_15(clock, reset, enable, direction, out_of_18_15, out_of_19_14, out_of_19_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_16(clock, reset, enable, direction, out_of_18_16, out_of_19_15, out_of_19_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_17(clock, reset, enable, direction, out_of_18_17, out_of_19_16, out_of_19_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_18(clock, reset, enable, direction, out_of_18_18, out_of_19_17, out_of_19_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_19(clock, reset, enable, direction, out_of_18_19, out_of_19_18, out_of_19_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_20(clock, reset, enable, direction, out_of_18_20, out_of_19_19, out_of_19_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_21(clock, reset, enable, direction, out_of_18_21, out_of_19_20, out_of_19_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_22(clock, reset, enable, direction, out_of_18_22, out_of_19_21, out_of_19_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_23(clock, reset, enable, direction, out_of_18_23, out_of_19_22, out_of_19_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_24(clock, reset, enable, direction, out_of_18_24, out_of_19_23, out_of_19_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_25(clock, reset, enable, direction, out_of_18_25, out_of_19_24, out_of_19_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_26(clock, reset, enable, direction, out_of_18_26, out_of_19_25, out_of_19_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_27(clock, reset, enable, direction, out_of_18_27, out_of_19_26, out_of_19_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_28(clock, reset, enable, direction, out_of_18_28, out_of_19_27, out_of_19_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_29(clock, reset, enable, direction, out_of_18_29, out_of_19_28, out_of_19_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_30(clock, reset, enable, direction, out_of_18_30, out_of_19_29, out_of_19_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_19_31(clock, reset, enable, direction, out_of_18_31, out_of_19_30, out_of_19_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_0(clock, reset, enable, direction, out_of_19_0, in_20, out_of_20_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_1(clock, reset, enable, direction, out_of_19_1, out_of_20_0, out_of_20_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_2(clock, reset, enable, direction, out_of_19_2, out_of_20_1, out_of_20_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_3(clock, reset, enable, direction, out_of_19_3, out_of_20_2, out_of_20_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_4(clock, reset, enable, direction, out_of_19_4, out_of_20_3, out_of_20_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_5(clock, reset, enable, direction, out_of_19_5, out_of_20_4, out_of_20_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_6(clock, reset, enable, direction, out_of_19_6, out_of_20_5, out_of_20_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_7(clock, reset, enable, direction, out_of_19_7, out_of_20_6, out_of_20_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_8(clock, reset, enable, direction, out_of_19_8, out_of_20_7, out_of_20_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_9(clock, reset, enable, direction, out_of_19_9, out_of_20_8, out_of_20_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_10(clock, reset, enable, direction, out_of_19_10, out_of_20_9, out_of_20_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_11(clock, reset, enable, direction, out_of_19_11, out_of_20_10, out_of_20_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_12(clock, reset, enable, direction, out_of_19_12, out_of_20_11, out_of_20_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_13(clock, reset, enable, direction, out_of_19_13, out_of_20_12, out_of_20_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_14(clock, reset, enable, direction, out_of_19_14, out_of_20_13, out_of_20_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_15(clock, reset, enable, direction, out_of_19_15, out_of_20_14, out_of_20_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_16(clock, reset, enable, direction, out_of_19_16, out_of_20_15, out_of_20_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_17(clock, reset, enable, direction, out_of_19_17, out_of_20_16, out_of_20_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_18(clock, reset, enable, direction, out_of_19_18, out_of_20_17, out_of_20_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_19(clock, reset, enable, direction, out_of_19_19, out_of_20_18, out_of_20_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_20(clock, reset, enable, direction, out_of_19_20, out_of_20_19, out_of_20_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_21(clock, reset, enable, direction, out_of_19_21, out_of_20_20, out_of_20_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_22(clock, reset, enable, direction, out_of_19_22, out_of_20_21, out_of_20_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_23(clock, reset, enable, direction, out_of_19_23, out_of_20_22, out_of_20_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_24(clock, reset, enable, direction, out_of_19_24, out_of_20_23, out_of_20_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_25(clock, reset, enable, direction, out_of_19_25, out_of_20_24, out_of_20_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_26(clock, reset, enable, direction, out_of_19_26, out_of_20_25, out_of_20_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_27(clock, reset, enable, direction, out_of_19_27, out_of_20_26, out_of_20_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_28(clock, reset, enable, direction, out_of_19_28, out_of_20_27, out_of_20_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_29(clock, reset, enable, direction, out_of_19_29, out_of_20_28, out_of_20_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_30(clock, reset, enable, direction, out_of_19_30, out_of_20_29, out_of_20_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_20_31(clock, reset, enable, direction, out_of_19_31, out_of_20_30, out_of_20_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_0(clock, reset, enable, direction, out_of_20_0, in_21, out_of_21_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_1(clock, reset, enable, direction, out_of_20_1, out_of_21_0, out_of_21_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_2(clock, reset, enable, direction, out_of_20_2, out_of_21_1, out_of_21_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_3(clock, reset, enable, direction, out_of_20_3, out_of_21_2, out_of_21_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_4(clock, reset, enable, direction, out_of_20_4, out_of_21_3, out_of_21_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_5(clock, reset, enable, direction, out_of_20_5, out_of_21_4, out_of_21_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_6(clock, reset, enable, direction, out_of_20_6, out_of_21_5, out_of_21_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_7(clock, reset, enable, direction, out_of_20_7, out_of_21_6, out_of_21_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_8(clock, reset, enable, direction, out_of_20_8, out_of_21_7, out_of_21_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_9(clock, reset, enable, direction, out_of_20_9, out_of_21_8, out_of_21_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_10(clock, reset, enable, direction, out_of_20_10, out_of_21_9, out_of_21_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_11(clock, reset, enable, direction, out_of_20_11, out_of_21_10, out_of_21_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_12(clock, reset, enable, direction, out_of_20_12, out_of_21_11, out_of_21_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_13(clock, reset, enable, direction, out_of_20_13, out_of_21_12, out_of_21_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_14(clock, reset, enable, direction, out_of_20_14, out_of_21_13, out_of_21_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_15(clock, reset, enable, direction, out_of_20_15, out_of_21_14, out_of_21_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_16(clock, reset, enable, direction, out_of_20_16, out_of_21_15, out_of_21_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_17(clock, reset, enable, direction, out_of_20_17, out_of_21_16, out_of_21_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_18(clock, reset, enable, direction, out_of_20_18, out_of_21_17, out_of_21_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_19(clock, reset, enable, direction, out_of_20_19, out_of_21_18, out_of_21_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_20(clock, reset, enable, direction, out_of_20_20, out_of_21_19, out_of_21_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_21(clock, reset, enable, direction, out_of_20_21, out_of_21_20, out_of_21_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_22(clock, reset, enable, direction, out_of_20_22, out_of_21_21, out_of_21_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_23(clock, reset, enable, direction, out_of_20_23, out_of_21_22, out_of_21_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_24(clock, reset, enable, direction, out_of_20_24, out_of_21_23, out_of_21_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_25(clock, reset, enable, direction, out_of_20_25, out_of_21_24, out_of_21_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_26(clock, reset, enable, direction, out_of_20_26, out_of_21_25, out_of_21_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_27(clock, reset, enable, direction, out_of_20_27, out_of_21_26, out_of_21_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_28(clock, reset, enable, direction, out_of_20_28, out_of_21_27, out_of_21_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_29(clock, reset, enable, direction, out_of_20_29, out_of_21_28, out_of_21_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_30(clock, reset, enable, direction, out_of_20_30, out_of_21_29, out_of_21_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_21_31(clock, reset, enable, direction, out_of_20_31, out_of_21_30, out_of_21_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_0(clock, reset, enable, direction, out_of_21_0, in_22, out_of_22_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_1(clock, reset, enable, direction, out_of_21_1, out_of_22_0, out_of_22_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_2(clock, reset, enable, direction, out_of_21_2, out_of_22_1, out_of_22_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_3(clock, reset, enable, direction, out_of_21_3, out_of_22_2, out_of_22_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_4(clock, reset, enable, direction, out_of_21_4, out_of_22_3, out_of_22_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_5(clock, reset, enable, direction, out_of_21_5, out_of_22_4, out_of_22_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_6(clock, reset, enable, direction, out_of_21_6, out_of_22_5, out_of_22_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_7(clock, reset, enable, direction, out_of_21_7, out_of_22_6, out_of_22_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_8(clock, reset, enable, direction, out_of_21_8, out_of_22_7, out_of_22_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_9(clock, reset, enable, direction, out_of_21_9, out_of_22_8, out_of_22_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_10(clock, reset, enable, direction, out_of_21_10, out_of_22_9, out_of_22_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_11(clock, reset, enable, direction, out_of_21_11, out_of_22_10, out_of_22_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_12(clock, reset, enable, direction, out_of_21_12, out_of_22_11, out_of_22_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_13(clock, reset, enable, direction, out_of_21_13, out_of_22_12, out_of_22_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_14(clock, reset, enable, direction, out_of_21_14, out_of_22_13, out_of_22_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_15(clock, reset, enable, direction, out_of_21_15, out_of_22_14, out_of_22_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_16(clock, reset, enable, direction, out_of_21_16, out_of_22_15, out_of_22_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_17(clock, reset, enable, direction, out_of_21_17, out_of_22_16, out_of_22_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_18(clock, reset, enable, direction, out_of_21_18, out_of_22_17, out_of_22_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_19(clock, reset, enable, direction, out_of_21_19, out_of_22_18, out_of_22_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_20(clock, reset, enable, direction, out_of_21_20, out_of_22_19, out_of_22_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_21(clock, reset, enable, direction, out_of_21_21, out_of_22_20, out_of_22_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_22(clock, reset, enable, direction, out_of_21_22, out_of_22_21, out_of_22_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_23(clock, reset, enable, direction, out_of_21_23, out_of_22_22, out_of_22_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_24(clock, reset, enable, direction, out_of_21_24, out_of_22_23, out_of_22_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_25(clock, reset, enable, direction, out_of_21_25, out_of_22_24, out_of_22_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_26(clock, reset, enable, direction, out_of_21_26, out_of_22_25, out_of_22_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_27(clock, reset, enable, direction, out_of_21_27, out_of_22_26, out_of_22_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_28(clock, reset, enable, direction, out_of_21_28, out_of_22_27, out_of_22_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_29(clock, reset, enable, direction, out_of_21_29, out_of_22_28, out_of_22_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_30(clock, reset, enable, direction, out_of_21_30, out_of_22_29, out_of_22_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_22_31(clock, reset, enable, direction, out_of_21_31, out_of_22_30, out_of_22_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_0(clock, reset, enable, direction, out_of_22_0, in_23, out_of_23_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_1(clock, reset, enable, direction, out_of_22_1, out_of_23_0, out_of_23_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_2(clock, reset, enable, direction, out_of_22_2, out_of_23_1, out_of_23_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_3(clock, reset, enable, direction, out_of_22_3, out_of_23_2, out_of_23_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_4(clock, reset, enable, direction, out_of_22_4, out_of_23_3, out_of_23_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_5(clock, reset, enable, direction, out_of_22_5, out_of_23_4, out_of_23_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_6(clock, reset, enable, direction, out_of_22_6, out_of_23_5, out_of_23_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_7(clock, reset, enable, direction, out_of_22_7, out_of_23_6, out_of_23_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_8(clock, reset, enable, direction, out_of_22_8, out_of_23_7, out_of_23_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_9(clock, reset, enable, direction, out_of_22_9, out_of_23_8, out_of_23_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_10(clock, reset, enable, direction, out_of_22_10, out_of_23_9, out_of_23_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_11(clock, reset, enable, direction, out_of_22_11, out_of_23_10, out_of_23_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_12(clock, reset, enable, direction, out_of_22_12, out_of_23_11, out_of_23_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_13(clock, reset, enable, direction, out_of_22_13, out_of_23_12, out_of_23_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_14(clock, reset, enable, direction, out_of_22_14, out_of_23_13, out_of_23_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_15(clock, reset, enable, direction, out_of_22_15, out_of_23_14, out_of_23_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_16(clock, reset, enable, direction, out_of_22_16, out_of_23_15, out_of_23_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_17(clock, reset, enable, direction, out_of_22_17, out_of_23_16, out_of_23_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_18(clock, reset, enable, direction, out_of_22_18, out_of_23_17, out_of_23_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_19(clock, reset, enable, direction, out_of_22_19, out_of_23_18, out_of_23_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_20(clock, reset, enable, direction, out_of_22_20, out_of_23_19, out_of_23_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_21(clock, reset, enable, direction, out_of_22_21, out_of_23_20, out_of_23_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_22(clock, reset, enable, direction, out_of_22_22, out_of_23_21, out_of_23_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_23(clock, reset, enable, direction, out_of_22_23, out_of_23_22, out_of_23_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_24(clock, reset, enable, direction, out_of_22_24, out_of_23_23, out_of_23_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_25(clock, reset, enable, direction, out_of_22_25, out_of_23_24, out_of_23_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_26(clock, reset, enable, direction, out_of_22_26, out_of_23_25, out_of_23_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_27(clock, reset, enable, direction, out_of_22_27, out_of_23_26, out_of_23_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_28(clock, reset, enable, direction, out_of_22_28, out_of_23_27, out_of_23_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_29(clock, reset, enable, direction, out_of_22_29, out_of_23_28, out_of_23_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_30(clock, reset, enable, direction, out_of_22_30, out_of_23_29, out_of_23_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_23_31(clock, reset, enable, direction, out_of_22_31, out_of_23_30, out_of_23_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_0(clock, reset, enable, direction, out_of_23_0, in_24, out_of_24_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_1(clock, reset, enable, direction, out_of_23_1, out_of_24_0, out_of_24_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_2(clock, reset, enable, direction, out_of_23_2, out_of_24_1, out_of_24_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_3(clock, reset, enable, direction, out_of_23_3, out_of_24_2, out_of_24_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_4(clock, reset, enable, direction, out_of_23_4, out_of_24_3, out_of_24_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_5(clock, reset, enable, direction, out_of_23_5, out_of_24_4, out_of_24_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_6(clock, reset, enable, direction, out_of_23_6, out_of_24_5, out_of_24_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_7(clock, reset, enable, direction, out_of_23_7, out_of_24_6, out_of_24_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_8(clock, reset, enable, direction, out_of_23_8, out_of_24_7, out_of_24_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_9(clock, reset, enable, direction, out_of_23_9, out_of_24_8, out_of_24_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_10(clock, reset, enable, direction, out_of_23_10, out_of_24_9, out_of_24_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_11(clock, reset, enable, direction, out_of_23_11, out_of_24_10, out_of_24_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_12(clock, reset, enable, direction, out_of_23_12, out_of_24_11, out_of_24_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_13(clock, reset, enable, direction, out_of_23_13, out_of_24_12, out_of_24_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_14(clock, reset, enable, direction, out_of_23_14, out_of_24_13, out_of_24_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_15(clock, reset, enable, direction, out_of_23_15, out_of_24_14, out_of_24_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_16(clock, reset, enable, direction, out_of_23_16, out_of_24_15, out_of_24_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_17(clock, reset, enable, direction, out_of_23_17, out_of_24_16, out_of_24_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_18(clock, reset, enable, direction, out_of_23_18, out_of_24_17, out_of_24_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_19(clock, reset, enable, direction, out_of_23_19, out_of_24_18, out_of_24_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_20(clock, reset, enable, direction, out_of_23_20, out_of_24_19, out_of_24_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_21(clock, reset, enable, direction, out_of_23_21, out_of_24_20, out_of_24_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_22(clock, reset, enable, direction, out_of_23_22, out_of_24_21, out_of_24_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_23(clock, reset, enable, direction, out_of_23_23, out_of_24_22, out_of_24_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_24(clock, reset, enable, direction, out_of_23_24, out_of_24_23, out_of_24_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_25(clock, reset, enable, direction, out_of_23_25, out_of_24_24, out_of_24_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_26(clock, reset, enable, direction, out_of_23_26, out_of_24_25, out_of_24_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_27(clock, reset, enable, direction, out_of_23_27, out_of_24_26, out_of_24_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_28(clock, reset, enable, direction, out_of_23_28, out_of_24_27, out_of_24_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_29(clock, reset, enable, direction, out_of_23_29, out_of_24_28, out_of_24_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_30(clock, reset, enable, direction, out_of_23_30, out_of_24_29, out_of_24_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_24_31(clock, reset, enable, direction, out_of_23_31, out_of_24_30, out_of_24_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_0(clock, reset, enable, direction, out_of_24_0, in_25, out_of_25_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_1(clock, reset, enable, direction, out_of_24_1, out_of_25_0, out_of_25_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_2(clock, reset, enable, direction, out_of_24_2, out_of_25_1, out_of_25_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_3(clock, reset, enable, direction, out_of_24_3, out_of_25_2, out_of_25_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_4(clock, reset, enable, direction, out_of_24_4, out_of_25_3, out_of_25_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_5(clock, reset, enable, direction, out_of_24_5, out_of_25_4, out_of_25_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_6(clock, reset, enable, direction, out_of_24_6, out_of_25_5, out_of_25_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_7(clock, reset, enable, direction, out_of_24_7, out_of_25_6, out_of_25_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_8(clock, reset, enable, direction, out_of_24_8, out_of_25_7, out_of_25_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_9(clock, reset, enable, direction, out_of_24_9, out_of_25_8, out_of_25_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_10(clock, reset, enable, direction, out_of_24_10, out_of_25_9, out_of_25_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_11(clock, reset, enable, direction, out_of_24_11, out_of_25_10, out_of_25_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_12(clock, reset, enable, direction, out_of_24_12, out_of_25_11, out_of_25_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_13(clock, reset, enable, direction, out_of_24_13, out_of_25_12, out_of_25_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_14(clock, reset, enable, direction, out_of_24_14, out_of_25_13, out_of_25_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_15(clock, reset, enable, direction, out_of_24_15, out_of_25_14, out_of_25_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_16(clock, reset, enable, direction, out_of_24_16, out_of_25_15, out_of_25_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_17(clock, reset, enable, direction, out_of_24_17, out_of_25_16, out_of_25_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_18(clock, reset, enable, direction, out_of_24_18, out_of_25_17, out_of_25_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_19(clock, reset, enable, direction, out_of_24_19, out_of_25_18, out_of_25_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_20(clock, reset, enable, direction, out_of_24_20, out_of_25_19, out_of_25_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_21(clock, reset, enable, direction, out_of_24_21, out_of_25_20, out_of_25_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_22(clock, reset, enable, direction, out_of_24_22, out_of_25_21, out_of_25_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_23(clock, reset, enable, direction, out_of_24_23, out_of_25_22, out_of_25_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_24(clock, reset, enable, direction, out_of_24_24, out_of_25_23, out_of_25_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_25(clock, reset, enable, direction, out_of_24_25, out_of_25_24, out_of_25_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_26(clock, reset, enable, direction, out_of_24_26, out_of_25_25, out_of_25_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_27(clock, reset, enable, direction, out_of_24_27, out_of_25_26, out_of_25_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_28(clock, reset, enable, direction, out_of_24_28, out_of_25_27, out_of_25_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_29(clock, reset, enable, direction, out_of_24_29, out_of_25_28, out_of_25_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_30(clock, reset, enable, direction, out_of_24_30, out_of_25_29, out_of_25_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_25_31(clock, reset, enable, direction, out_of_24_31, out_of_25_30, out_of_25_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_0(clock, reset, enable, direction, out_of_25_0, in_26, out_of_26_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_1(clock, reset, enable, direction, out_of_25_1, out_of_26_0, out_of_26_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_2(clock, reset, enable, direction, out_of_25_2, out_of_26_1, out_of_26_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_3(clock, reset, enable, direction, out_of_25_3, out_of_26_2, out_of_26_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_4(clock, reset, enable, direction, out_of_25_4, out_of_26_3, out_of_26_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_5(clock, reset, enable, direction, out_of_25_5, out_of_26_4, out_of_26_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_6(clock, reset, enable, direction, out_of_25_6, out_of_26_5, out_of_26_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_7(clock, reset, enable, direction, out_of_25_7, out_of_26_6, out_of_26_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_8(clock, reset, enable, direction, out_of_25_8, out_of_26_7, out_of_26_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_9(clock, reset, enable, direction, out_of_25_9, out_of_26_8, out_of_26_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_10(clock, reset, enable, direction, out_of_25_10, out_of_26_9, out_of_26_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_11(clock, reset, enable, direction, out_of_25_11, out_of_26_10, out_of_26_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_12(clock, reset, enable, direction, out_of_25_12, out_of_26_11, out_of_26_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_13(clock, reset, enable, direction, out_of_25_13, out_of_26_12, out_of_26_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_14(clock, reset, enable, direction, out_of_25_14, out_of_26_13, out_of_26_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_15(clock, reset, enable, direction, out_of_25_15, out_of_26_14, out_of_26_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_16(clock, reset, enable, direction, out_of_25_16, out_of_26_15, out_of_26_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_17(clock, reset, enable, direction, out_of_25_17, out_of_26_16, out_of_26_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_18(clock, reset, enable, direction, out_of_25_18, out_of_26_17, out_of_26_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_19(clock, reset, enable, direction, out_of_25_19, out_of_26_18, out_of_26_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_20(clock, reset, enable, direction, out_of_25_20, out_of_26_19, out_of_26_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_21(clock, reset, enable, direction, out_of_25_21, out_of_26_20, out_of_26_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_22(clock, reset, enable, direction, out_of_25_22, out_of_26_21, out_of_26_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_23(clock, reset, enable, direction, out_of_25_23, out_of_26_22, out_of_26_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_24(clock, reset, enable, direction, out_of_25_24, out_of_26_23, out_of_26_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_25(clock, reset, enable, direction, out_of_25_25, out_of_26_24, out_of_26_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_26(clock, reset, enable, direction, out_of_25_26, out_of_26_25, out_of_26_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_27(clock, reset, enable, direction, out_of_25_27, out_of_26_26, out_of_26_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_28(clock, reset, enable, direction, out_of_25_28, out_of_26_27, out_of_26_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_29(clock, reset, enable, direction, out_of_25_29, out_of_26_28, out_of_26_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_30(clock, reset, enable, direction, out_of_25_30, out_of_26_29, out_of_26_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_26_31(clock, reset, enable, direction, out_of_25_31, out_of_26_30, out_of_26_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_0(clock, reset, enable, direction, out_of_26_0, in_27, out_of_27_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_1(clock, reset, enable, direction, out_of_26_1, out_of_27_0, out_of_27_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_2(clock, reset, enable, direction, out_of_26_2, out_of_27_1, out_of_27_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_3(clock, reset, enable, direction, out_of_26_3, out_of_27_2, out_of_27_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_4(clock, reset, enable, direction, out_of_26_4, out_of_27_3, out_of_27_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_5(clock, reset, enable, direction, out_of_26_5, out_of_27_4, out_of_27_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_6(clock, reset, enable, direction, out_of_26_6, out_of_27_5, out_of_27_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_7(clock, reset, enable, direction, out_of_26_7, out_of_27_6, out_of_27_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_8(clock, reset, enable, direction, out_of_26_8, out_of_27_7, out_of_27_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_9(clock, reset, enable, direction, out_of_26_9, out_of_27_8, out_of_27_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_10(clock, reset, enable, direction, out_of_26_10, out_of_27_9, out_of_27_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_11(clock, reset, enable, direction, out_of_26_11, out_of_27_10, out_of_27_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_12(clock, reset, enable, direction, out_of_26_12, out_of_27_11, out_of_27_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_13(clock, reset, enable, direction, out_of_26_13, out_of_27_12, out_of_27_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_14(clock, reset, enable, direction, out_of_26_14, out_of_27_13, out_of_27_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_15(clock, reset, enable, direction, out_of_26_15, out_of_27_14, out_of_27_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_16(clock, reset, enable, direction, out_of_26_16, out_of_27_15, out_of_27_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_17(clock, reset, enable, direction, out_of_26_17, out_of_27_16, out_of_27_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_18(clock, reset, enable, direction, out_of_26_18, out_of_27_17, out_of_27_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_19(clock, reset, enable, direction, out_of_26_19, out_of_27_18, out_of_27_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_20(clock, reset, enable, direction, out_of_26_20, out_of_27_19, out_of_27_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_21(clock, reset, enable, direction, out_of_26_21, out_of_27_20, out_of_27_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_22(clock, reset, enable, direction, out_of_26_22, out_of_27_21, out_of_27_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_23(clock, reset, enable, direction, out_of_26_23, out_of_27_22, out_of_27_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_24(clock, reset, enable, direction, out_of_26_24, out_of_27_23, out_of_27_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_25(clock, reset, enable, direction, out_of_26_25, out_of_27_24, out_of_27_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_26(clock, reset, enable, direction, out_of_26_26, out_of_27_25, out_of_27_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_27(clock, reset, enable, direction, out_of_26_27, out_of_27_26, out_of_27_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_28(clock, reset, enable, direction, out_of_26_28, out_of_27_27, out_of_27_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_29(clock, reset, enable, direction, out_of_26_29, out_of_27_28, out_of_27_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_30(clock, reset, enable, direction, out_of_26_30, out_of_27_29, out_of_27_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_27_31(clock, reset, enable, direction, out_of_26_31, out_of_27_30, out_of_27_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_0(clock, reset, enable, direction, out_of_27_0, in_28, out_of_28_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_1(clock, reset, enable, direction, out_of_27_1, out_of_28_0, out_of_28_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_2(clock, reset, enable, direction, out_of_27_2, out_of_28_1, out_of_28_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_3(clock, reset, enable, direction, out_of_27_3, out_of_28_2, out_of_28_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_4(clock, reset, enable, direction, out_of_27_4, out_of_28_3, out_of_28_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_5(clock, reset, enable, direction, out_of_27_5, out_of_28_4, out_of_28_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_6(clock, reset, enable, direction, out_of_27_6, out_of_28_5, out_of_28_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_7(clock, reset, enable, direction, out_of_27_7, out_of_28_6, out_of_28_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_8(clock, reset, enable, direction, out_of_27_8, out_of_28_7, out_of_28_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_9(clock, reset, enable, direction, out_of_27_9, out_of_28_8, out_of_28_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_10(clock, reset, enable, direction, out_of_27_10, out_of_28_9, out_of_28_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_11(clock, reset, enable, direction, out_of_27_11, out_of_28_10, out_of_28_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_12(clock, reset, enable, direction, out_of_27_12, out_of_28_11, out_of_28_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_13(clock, reset, enable, direction, out_of_27_13, out_of_28_12, out_of_28_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_14(clock, reset, enable, direction, out_of_27_14, out_of_28_13, out_of_28_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_15(clock, reset, enable, direction, out_of_27_15, out_of_28_14, out_of_28_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_16(clock, reset, enable, direction, out_of_27_16, out_of_28_15, out_of_28_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_17(clock, reset, enable, direction, out_of_27_17, out_of_28_16, out_of_28_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_18(clock, reset, enable, direction, out_of_27_18, out_of_28_17, out_of_28_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_19(clock, reset, enable, direction, out_of_27_19, out_of_28_18, out_of_28_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_20(clock, reset, enable, direction, out_of_27_20, out_of_28_19, out_of_28_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_21(clock, reset, enable, direction, out_of_27_21, out_of_28_20, out_of_28_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_22(clock, reset, enable, direction, out_of_27_22, out_of_28_21, out_of_28_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_23(clock, reset, enable, direction, out_of_27_23, out_of_28_22, out_of_28_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_24(clock, reset, enable, direction, out_of_27_24, out_of_28_23, out_of_28_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_25(clock, reset, enable, direction, out_of_27_25, out_of_28_24, out_of_28_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_26(clock, reset, enable, direction, out_of_27_26, out_of_28_25, out_of_28_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_27(clock, reset, enable, direction, out_of_27_27, out_of_28_26, out_of_28_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_28(clock, reset, enable, direction, out_of_27_28, out_of_28_27, out_of_28_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_29(clock, reset, enable, direction, out_of_27_29, out_of_28_28, out_of_28_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_30(clock, reset, enable, direction, out_of_27_30, out_of_28_29, out_of_28_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_28_31(clock, reset, enable, direction, out_of_27_31, out_of_28_30, out_of_28_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_0(clock, reset, enable, direction, out_of_28_0, in_29, out_of_29_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_1(clock, reset, enable, direction, out_of_28_1, out_of_29_0, out_of_29_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_2(clock, reset, enable, direction, out_of_28_2, out_of_29_1, out_of_29_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_3(clock, reset, enable, direction, out_of_28_3, out_of_29_2, out_of_29_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_4(clock, reset, enable, direction, out_of_28_4, out_of_29_3, out_of_29_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_5(clock, reset, enable, direction, out_of_28_5, out_of_29_4, out_of_29_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_6(clock, reset, enable, direction, out_of_28_6, out_of_29_5, out_of_29_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_7(clock, reset, enable, direction, out_of_28_7, out_of_29_6, out_of_29_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_8(clock, reset, enable, direction, out_of_28_8, out_of_29_7, out_of_29_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_9(clock, reset, enable, direction, out_of_28_9, out_of_29_8, out_of_29_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_10(clock, reset, enable, direction, out_of_28_10, out_of_29_9, out_of_29_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_11(clock, reset, enable, direction, out_of_28_11, out_of_29_10, out_of_29_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_12(clock, reset, enable, direction, out_of_28_12, out_of_29_11, out_of_29_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_13(clock, reset, enable, direction, out_of_28_13, out_of_29_12, out_of_29_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_14(clock, reset, enable, direction, out_of_28_14, out_of_29_13, out_of_29_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_15(clock, reset, enable, direction, out_of_28_15, out_of_29_14, out_of_29_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_16(clock, reset, enable, direction, out_of_28_16, out_of_29_15, out_of_29_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_17(clock, reset, enable, direction, out_of_28_17, out_of_29_16, out_of_29_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_18(clock, reset, enable, direction, out_of_28_18, out_of_29_17, out_of_29_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_19(clock, reset, enable, direction, out_of_28_19, out_of_29_18, out_of_29_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_20(clock, reset, enable, direction, out_of_28_20, out_of_29_19, out_of_29_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_21(clock, reset, enable, direction, out_of_28_21, out_of_29_20, out_of_29_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_22(clock, reset, enable, direction, out_of_28_22, out_of_29_21, out_of_29_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_23(clock, reset, enable, direction, out_of_28_23, out_of_29_22, out_of_29_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_24(clock, reset, enable, direction, out_of_28_24, out_of_29_23, out_of_29_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_25(clock, reset, enable, direction, out_of_28_25, out_of_29_24, out_of_29_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_26(clock, reset, enable, direction, out_of_28_26, out_of_29_25, out_of_29_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_27(clock, reset, enable, direction, out_of_28_27, out_of_29_26, out_of_29_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_28(clock, reset, enable, direction, out_of_28_28, out_of_29_27, out_of_29_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_29(clock, reset, enable, direction, out_of_28_29, out_of_29_28, out_of_29_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_30(clock, reset, enable, direction, out_of_28_30, out_of_29_29, out_of_29_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_29_31(clock, reset, enable, direction, out_of_28_31, out_of_29_30, out_of_29_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_0(clock, reset, enable, direction, out_of_29_0, in_30, out_of_30_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_1(clock, reset, enable, direction, out_of_29_1, out_of_30_0, out_of_30_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_2(clock, reset, enable, direction, out_of_29_2, out_of_30_1, out_of_30_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_3(clock, reset, enable, direction, out_of_29_3, out_of_30_2, out_of_30_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_4(clock, reset, enable, direction, out_of_29_4, out_of_30_3, out_of_30_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_5(clock, reset, enable, direction, out_of_29_5, out_of_30_4, out_of_30_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_6(clock, reset, enable, direction, out_of_29_6, out_of_30_5, out_of_30_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_7(clock, reset, enable, direction, out_of_29_7, out_of_30_6, out_of_30_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_8(clock, reset, enable, direction, out_of_29_8, out_of_30_7, out_of_30_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_9(clock, reset, enable, direction, out_of_29_9, out_of_30_8, out_of_30_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_10(clock, reset, enable, direction, out_of_29_10, out_of_30_9, out_of_30_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_11(clock, reset, enable, direction, out_of_29_11, out_of_30_10, out_of_30_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_12(clock, reset, enable, direction, out_of_29_12, out_of_30_11, out_of_30_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_13(clock, reset, enable, direction, out_of_29_13, out_of_30_12, out_of_30_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_14(clock, reset, enable, direction, out_of_29_14, out_of_30_13, out_of_30_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_15(clock, reset, enable, direction, out_of_29_15, out_of_30_14, out_of_30_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_16(clock, reset, enable, direction, out_of_29_16, out_of_30_15, out_of_30_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_17(clock, reset, enable, direction, out_of_29_17, out_of_30_16, out_of_30_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_18(clock, reset, enable, direction, out_of_29_18, out_of_30_17, out_of_30_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_19(clock, reset, enable, direction, out_of_29_19, out_of_30_18, out_of_30_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_20(clock, reset, enable, direction, out_of_29_20, out_of_30_19, out_of_30_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_21(clock, reset, enable, direction, out_of_29_21, out_of_30_20, out_of_30_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_22(clock, reset, enable, direction, out_of_29_22, out_of_30_21, out_of_30_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_23(clock, reset, enable, direction, out_of_29_23, out_of_30_22, out_of_30_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_24(clock, reset, enable, direction, out_of_29_24, out_of_30_23, out_of_30_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_25(clock, reset, enable, direction, out_of_29_25, out_of_30_24, out_of_30_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_26(clock, reset, enable, direction, out_of_29_26, out_of_30_25, out_of_30_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_27(clock, reset, enable, direction, out_of_29_27, out_of_30_26, out_of_30_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_28(clock, reset, enable, direction, out_of_29_28, out_of_30_27, out_of_30_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_29(clock, reset, enable, direction, out_of_29_29, out_of_30_28, out_of_30_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_30(clock, reset, enable, direction, out_of_29_30, out_of_30_29, out_of_30_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_30_31(clock, reset, enable, direction, out_of_29_31, out_of_30_30, out_of_30_31);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_0(clock, reset, enable, direction, out_of_30_0, in_31, out_of_31_0);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_1(clock, reset, enable, direction, out_of_30_1, out_of_31_0, out_of_31_1);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_2(clock, reset, enable, direction, out_of_30_2, out_of_31_1, out_of_31_2);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_3(clock, reset, enable, direction, out_of_30_3, out_of_31_2, out_of_31_3);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_4(clock, reset, enable, direction, out_of_30_4, out_of_31_3, out_of_31_4);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_5(clock, reset, enable, direction, out_of_30_5, out_of_31_4, out_of_31_5);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_6(clock, reset, enable, direction, out_of_30_6, out_of_31_5, out_of_31_6);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_7(clock, reset, enable, direction, out_of_30_7, out_of_31_6, out_of_31_7);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_8(clock, reset, enable, direction, out_of_30_8, out_of_31_7, out_of_31_8);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_9(clock, reset, enable, direction, out_of_30_9, out_of_31_8, out_of_31_9);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_10(clock, reset, enable, direction, out_of_30_10, out_of_31_9, out_of_31_10);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_11(clock, reset, enable, direction, out_of_30_11, out_of_31_10, out_of_31_11);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_12(clock, reset, enable, direction, out_of_30_12, out_of_31_11, out_of_31_12);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_13(clock, reset, enable, direction, out_of_30_13, out_of_31_12, out_of_31_13);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_14(clock, reset, enable, direction, out_of_30_14, out_of_31_13, out_of_31_14);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_15(clock, reset, enable, direction, out_of_30_15, out_of_31_14, out_of_31_15);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_16(clock, reset, enable, direction, out_of_30_16, out_of_31_15, out_of_31_16);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_17(clock, reset, enable, direction, out_of_30_17, out_of_31_16, out_of_31_17);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_18(clock, reset, enable, direction, out_of_30_18, out_of_31_17, out_of_31_18);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_19(clock, reset, enable, direction, out_of_30_19, out_of_31_18, out_of_31_19);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_20(clock, reset, enable, direction, out_of_30_20, out_of_31_19, out_of_31_20);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_21(clock, reset, enable, direction, out_of_30_21, out_of_31_20, out_of_31_21);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_22(clock, reset, enable, direction, out_of_30_22, out_of_31_21, out_of_31_22);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_23(clock, reset, enable, direction, out_of_30_23, out_of_31_22, out_of_31_23);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_24(clock, reset, enable, direction, out_of_30_24, out_of_31_23, out_of_31_24);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_25(clock, reset, enable, direction, out_of_30_25, out_of_31_24, out_of_31_25);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_26(clock, reset, enable, direction, out_of_30_26, out_of_31_25, out_of_31_26);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_27(clock, reset, enable, direction, out_of_30_27, out_of_31_26, out_of_31_27);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_28(clock, reset, enable, direction, out_of_30_28, out_of_31_27, out_of_31_28);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_29(clock, reset, enable, direction, out_of_30_29, out_of_31_28, out_of_31_29);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_30(clock, reset, enable, direction, out_of_30_30, out_of_31_29, out_of_31_30);
transpose_buffer_cell #(DATA_WIDTH) tb_cell_31_31(clock, reset, enable, direction, out_of_30_31, out_of_31_30, out_of_31_31);

assign out_0  = (direction) ? out_of_0_31  : out_of_31_31;
assign out_1  = (direction) ? out_of_1_31  : out_of_31_30;
assign out_2  = (direction) ? out_of_2_31  : out_of_31_29;
assign out_3  = (direction) ? out_of_3_31  : out_of_31_28;
assign out_4  = (direction) ? out_of_4_31  : out_of_31_27;
assign out_5  = (direction) ? out_of_5_31  : out_of_31_26;
assign out_6  = (direction) ? out_of_6_31  : out_of_31_25;
assign out_7  = (direction) ? out_of_7_31  : out_of_31_24;
assign out_8  = (direction) ? out_of_8_31  : out_of_31_23;
assign out_9  = (direction) ? out_of_9_31  : out_of_31_22;
assign out_10 = (direction) ? out_of_10_31 : out_of_31_21;
assign out_11 = (direction) ? out_of_11_31 : out_of_31_20;
assign out_12 = (direction) ? out_of_12_31 : out_of_31_19;
assign out_13 = (direction) ? out_of_13_31 : out_of_31_18;
assign out_14 = (direction) ? out_of_14_31 : out_of_31_17;
assign out_15 = (direction) ? out_of_15_31 : out_of_31_16;
assign out_16 = (direction) ? out_of_16_31 : out_of_31_15;
assign out_17 = (direction) ? out_of_17_31 : out_of_31_14;
assign out_18 = (direction) ? out_of_18_31 : out_of_31_13;
assign out_19 = (direction) ? out_of_19_31 : out_of_31_12;
assign out_20 = (direction) ? out_of_20_31 : out_of_31_11;
assign out_21 = (direction) ? out_of_21_31 : out_of_31_10;
assign out_22 = (direction) ? out_of_22_31 : out_of_31_9 ;
assign out_23 = (direction) ? out_of_23_31 : out_of_31_8 ;
assign out_24 = (direction) ? out_of_24_31 : out_of_31_7 ;
assign out_25 = (direction) ? out_of_25_31 : out_of_31_6 ;
assign out_26 = (direction) ? out_of_26_31 : out_of_31_5 ;
assign out_27 = (direction) ? out_of_27_31 : out_of_31_4 ;
assign out_28 = (direction) ? out_of_28_31 : out_of_31_3 ;
assign out_29 = (direction) ? out_of_29_31 : out_of_31_2 ;
assign out_30 = (direction) ? out_of_30_31 : out_of_31_1 ;
assign out_31 = (direction) ? out_of_31_31 : out_of_31_0 ;

endmodule
