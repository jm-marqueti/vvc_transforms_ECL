module dct2_32 (input signed [15:0]X[0:31], 
output signed [16:0]Ye[0:15],
output signed [26:0]Yo[0:15]); 


//even-odd decomp
wire signed [16:0] E[0:15], O[0:15];

generate
genvar i;
	for (i = 0; i < 16; i = i + 1) begin: dcmploop
		decomp_0 decomposicao(X[i], X[31-i], E[i], O[i]);
	end
endgenerate


	//EVEN

assign Ye = E;

	//ODD (T2O)
	
wire signed [26:0] x4[0:15], x13[0:15], x22[0:15], x31[0:15],x38[0:15],x46[0:15],x54[0:15],x61[0:15],x67[0:15],x73[0:15],x78[0:15],x82[0:15],x85[0:15],x88[0:15],x90[0:15];

generate // SAU Setup
genvar j;
	for (j = 0; j < 16; j = j + 1) begin: oddSAUloop
		sau_16o sau_odd(O[j],x4[j], x13[j], x22[j], x31[j],x38[j],x46[j],x54[j],x61[j],x67[j],x73[j],x78[j],x82[j],x85[j],x88[j],x90[j]);
	end
endgenerate

			//Adder Trees
			
assign Yo[0]  = x90[0] + x90[1] + x88[2] + x85[3] + x82[4] + x78[5] + x73[6] + x67[7] + x61[8] + x54[9] + x46[10] + x38[11] + x31[12] + x22[13] + x13[14] +  x4[15];
assign Yo[1]  = x90[0] + x82[1] + x67[2] + x46[3] + x22[4] -  x4[5] - x31[6] - x54[7] - x73[8] - x85[9] - x90[10] - x88[11] - x78[12] - x61[13] - x38[14] - x13[15];
assign Yo[2]  = x88[0] + x67[1] + x31[2] - x13[3] - x54[4] - x82[5] - x90[6] - x78[7] - x46[8] -  x4[9] + x38[10] + x73[11] + x90[12] + x85[13] + x61[14] + x22[15];
assign Yo[3]  = x85[0] + x46[1] - x13[2] - x67[3] - x90[4] - x73[5] - x22[6] + x38[7] + x82[8] + x88[9] + x54[10] -  x4[11] - x61[12] - x90[13] - x78[14] - x31[15];
assign Yo[4]  = x82[0] + x22[1] - x54[2] - x90[3] - x61[4] + x13[5] + x78[6] + x85[7] + x31[8] - x46[9] - x90[10] - x67[11] +  x4[12] + x73[13] + x88[14] + x38[15];
assign Yo[5]  = x78[0] -  x4[1] - x82[2] - x73[3] + x13[4] + x85[5] + x67[6] - x22[7] - x88[8] - x61[9] + x31[10] + x90[11] + x54[12] - x38[13] - x90[14] - x46[15];
assign Yo[6]  = x73[0] - x31[1] - x90[2] - x22[3] + x78[4] + x67[5] - x38[6] - x90[7] - x13[8] + x82[9] + x61[10] - x46[11] - x88[12] -  x4[13] + x85[14] + x54[15];
assign Yo[7]  = x67[0] - x54[1] - x78[2] + x38[3] + x85[4] - x22[5] - x90[6] +  x4[7] + x90[8] + x13[9] - x88[10] - x31[11] + x82[12] + x46[13] - x73[14] - x61[15];
assign Yo[8]  = x61[0] - x73[1] - x46[2] + x82[3] + x31[4] - x88[5] - x13[6] + x90[7] -  x4[8] - x90[9] + x22[10] + x85[11] - x38[12] - x78[13] + x54[14] + x67[15];
assign Yo[9]  = x54[0] - x85[1] -  x4[2] + x88[3] - x46[4] - x61[5] + x82[6] + x13[7] - x90[8] + x38[9] + x67[10] - x78[11] - x22[12] + x90[13] - x31[14] - x73[15];
assign Yo[10] = x46[0] - x90[1] + x38[2] + x54[3] - x90[4] + x31[5] + x61[6] - x88[7] + x22[8] + x67[9] - x85[10] + x13[11] + x73[12] - x82[13] +  x4[14] + x78[15];
assign Yo[11] = x38[0] - x88[1] + x73[2] -  x4[3] - x67[4] + x90[5] - x46[6] - x31[7] + x85[8] - x78[9] + x13[10] + x61[11] - x90[12] + x54[13] + x22[14] - x82[15];
assign Yo[12] = x31[0] - x78[1] + x90[2] - x61[3] +  x4[4] + x54[5] - x88[6] + x82[7] - x38[8] - x22[9] + x73[10] - x90[11] + x67[12] - x13[13] - x46[14] + x85[15];
assign Yo[13] = x22[0] - x61[1] + x85[2] - x90[3] + x73[4] - x38[5] -  x4[6] + x46[7] - x78[8] + x90[9] - x82[10] + x54[11] - x13[12] - x31[13] + x67[14] - x88[15];
assign Yo[14] = x13[0] - x38[1] + x61[2] - x78[3] + x88[4] - x90[5] + x85[6] - x73[7] + x54[8] - x31[9] +  x4[10] + x22[11] - x46[12] + x67[13] - x82[14] + x90[15];
assign Yo[15] =  x4[0] - x13[1] + x22[2] - x31[3] + x38[4] - x46[5] + x54[6] - x61[7] + x67[8] - x73[9] + x78[10] - x82[11] + x85[12] - x88[13] + x90[14] - x90[15];


endmodule