module dst7_16(
input signed [8:0]X[15:0],
output signed [15:0]Y[15:0]);


// SAU

/*
// Adder Trees
assign Y[0] = x4[0] + x8[1] + x13[2] + x17[3] + x20[4] + x24[5] + x28[6] + x31[7] + x34[8] + x36[9] + x39[10] + x41[11] + x42[12] + x43[13] + x44[14] + x45[15];
assign Y[1] = x13[0] + x24[1] + x34[2] + x41[3] + x44[4] + x44[5] + x41[6] + x34[7] + x24[8] + x13[9] - x13[11] - x24[12] - x34[13] - x41[14] - x44[15];
assign Y[2] = x20[0] + x36[1] + x44[2] + x42[3] + x31[4] + x13[5] - x8[6] - x28[7] - x41[8] - x45[9] - x39[10] - x24[11] - x4[12] + x17[13] + x34[14] + x43[15];
assign Y[3] = x28[0] + x43[1] + x41[2] + x20[3] - x8[4] - x34[5] - x45[6] - x36[7] - x13[8] + x17[9] + x39[10] + x44[11] + x31[12] + x4[13] - x24[14] - x42[15];
assign Y[4] = x34[0] + x44[1] + x24[2] - x13[3] - x41[4] - x41[5] - x13[6] + x24[7] + x44[8] + x34[9] - x34[11] - x44[12] - x24[13] + x13[14] + x41[15];
assign Y[5] = x39[0] + x39[1] - x39[3] - x39[4] + x39[6] + x39[7] - x39[9] - x39[10] + x39[12] + x39[13] - x39[15];
assign Y[6] = x42[0] + x28[1] - x24[2] - x43[3] - x4[4] + x41[5] + x31[6] - x20[7] - x44[8] - x8[9] + x39[10] + x34[11] - x17[12] - x45[13] - x13[14] + x36[15];
assign Y[7] = x44[0] + x13[1] - x41[2] - x24[3] + x34[4] + x34[5] - x24[6] - x41[7] + x13[8] + x44[9] - x44[11] - x13[12] + x41[13] + x24[14] - x34[15];
assign Y[8] = x45[0] - x4[1] - x44[2] + x8[3] + x43[4] - x13[5] - x42[6] + x17[7] + x41[8] - x20[9] - x39[10] + x24[11] + x36[12] - x28[13] - x34[14] + x31[15];
assign Y[9] = x43[0] - x20[1] - x34[2] + x36[3] + x17[4] - x44[5] + x4[6] + x42[7] - x24[8] - x31[9] + x39[10] + x13[11] - x45[12] + x8[13] + x41[14] - x28[15];
assign Y[10] = x41[0] - x34[1] - x13[2] + x44[3] - x24[4] - x24[5] + x44[6] - x13[7] - x34[8] + x41[9] - x41[11] + x34[12] + x13[13] - x44[14] + x24[15];
assign Y[11] = x36[0] - x42[1] + x13[2] + x28[3] - x45[4] + x24[5] + x17[6] - x43[7] + x34[8] + x4[9] - x39[10] + x41[11] - x8[12] - x31[13] + x44[14] - x20[15];
assign Y[12] = x31[0] - x45[1] + x34[2] - x4[3] - x28[4] + x44[5] - x36[6] + x8[7] + x24[8] - x43[9] + x39[10] - x13[11] - x20[12] + x42[13] - x41[14] + x17[15];
assign Y[13] = x24[0] - x41[1] + x44[2] - x34[3] + x13[4] + x13[5] - x34[6] + x44[7] - x41[8] + x24[9] - x24[11] + x41[12] - x44[13] + x34[14] - x13[15];
assign Y[14] = x17[0] - x31[1] + x41[2] - x45[3] + x42[4] - x34[5] + x20[6] - x4[7] - x13[8] + x28[9] - x39[10] + x44[11] - x43[12] + x36[13] - x24[14] + x8[15];
assign Y[15] = x8[0] - x17[1] + x24[2] - x31[3] + x36[4] - x41[5] + x43[6] - x45[7] + x44[8] - x42[9] + x39[10] - x34[11] + x28[12] - x20[13] + x13[14] - x4[15];

*/
endmodule